<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="400" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-goa1.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.87322954,5.7016703,444)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-7">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9-2" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9-2" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6-2" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="386.56996" ns1:cy="46.494543" ns1:document-units="px" ns1:current-layer="g6112" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="5120" ns1:window-height="1376" ns1:window-x="0" ns1:window-y="27" ns1:window-maximized="1" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid15026"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-1092.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="639" x="-16" y="872.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-640)">
    <ns0:g id="g5895" transform="matrix(1.6596824,0,0,1.5988696,-623.10583,837.19119)">
      <ns0:g transform="matrix(0.29958781,0,0,0.29170899,321.78845,-7.042621)" id="g5467">
        <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:12.45934677;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 464.46875,123.03125 0,0.125 c -0.44393,-0.0201 -0.89409,-0.0194 -1.3125,-0.0312 -0.0201,-5e-4 -0.0415,-6e-5 -0.0625,0 l 0,-0.0312 c -35.47303,0 -52.12084,18.17885 -58.53125,35.53125 -4.16563,11.27597 -2.56542,24.58143 -0.90625,38.0625 0.61719,5.01479 1.38934,10.3782 2.25,15.90625 0.0523,1.53427 0.0953,3.02176 0.0625,4.25 -0.48198,18.0321 -6.73844,40.14561 -6.375,53.75 0.67291,25.18859 14.15792,41.81557 32.09375,50.3125 0.28216,0.13367 0.55942,0.27661 0.84375,0.40625 20.53214,9.97483 44.84145,10.69846 64.53125,-2 17.00609,-9.04566 29.375,-25.39691 29.375,-48.71875 0,-13.60924 -5.89302,-35.7179 -6.375,-53.75 -0.19564,-7.31935 1.4375,-21.90625 1.4375,-21.90625 1.53635,-7.2428 2.64168,-15.026 2.34375,-22.59375 -0.004,-0.10339 0.005,-0.20919 0,-0.3125 -0.11179,-3.85613 -0.64084,-7.56265 -1.6875,-11.03125 -0.11795,-0.39089 -0.24268,-0.77221 -0.375,-1.15625 -0.10094,-0.32527 -0.172,-0.64602 -0.28125,-0.96875 -0.60655,-1.79171 -1.42373,-3.60933 -2.375,-5.40625 -0.0677,-0.13829 -0.15051,-0.26913 -0.21875,-0.40625 C 507.06524,129.26972 486.89808,123.03135 464.46875,123.03135 Z" id="use3906-7-3"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="ccsccscsc" ns1:connector-curvature="0" id="path3896-9" d="m 471.25496,79.200587 5.30654,-28.587308 c 0.64849,-3.57802 1.26981,-7.661014 0.0259,-10.803791 -3.14471,-7.945086 -9.05873,-9.963605 -15.689,-9.963605 l -0.37971,0.0146 c -9.79602,0 -14.39338,5.126277 -16.16364,10.019502 l -3e-5,1e-6 c -1.15035,3.179726 -0.70845,6.93175 -0.25026,10.733293 0.74423,6.174786 2.22673,14.066104 3.59775,20.732961" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.30693826;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5509" d="m 460.5,28.862183 0,23" style="fill:none;stroke:#000000;stroke-width:0.30693826;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none"/>
      <ns0:rect ry="1.0234503" rx="0.90486509" y="35.253452" x="458.65408" height="11.488176" width="3.691813" id="rect5511" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:0.6138764;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 444,54.362183 c 5.14462,-1.307176 9.93443,-2.504355 16.4928,-2.499994 6.55838,-0.0044 11.34819,1.192829 16.49281,2.500005" style="fill:none;stroke:#000000;stroke-width:0.30693826;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" id="path5509-2-7"/>
    </ns0:g>
    <ns0:g transform="matrix(-1.4230531,0,0,1.4230531,588.13412,373.47398)" id="g3938">
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" id="rect3201" d="m 146.93753,371.19797 0,-129.07529 143.35232,0" style="color:#000000;fill:#000000;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:2.10814333;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 148.37105,270.089 c 0,-3.56432 2.88813,-6.45377 6.45085,-6.45377 l 156.25403,0" style="fill:none;stroke:#000000;stroke-width:0.70271444px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" id="path3995"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 146.93753,270.089 c 0,-3.56432 2.88813,-6.45377 6.45085,-6.45377 l 82.9074,0" style="fill:none;stroke:#000000;stroke-width:2.10814333;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" id="path3995-8"/>
      <ns0:g transform="matrix(-1.4335232,0,0,1.4341698,208.82881,250.97122)" ns1:label="#g5607" id="default-pointer-c-1" style="display:inline">
        <ns0:path style="color:#000000;fill:url(#linearGradient4726-2-9);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.49009043;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 Z" id="path5565-2" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path ns2:nodetypes="cccccccc" id="path6242-4" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 Z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.49009043;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="ccccccccccc" ns1:connector-curvature="0" id="rect12572-5" d="m 251.22895,340.05538 -17.67947,-18.16056 m -21.57129,-22.15829 -4.48672,-4.60881 7.09558,-7.09879 -26.35501,-2.02823 2.02732,26.3669 7.09558,-7.09878 10.99783,11.00279 m 10.93061,10.93554 33.27093,33.28595" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.70271444;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0.95;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:g transform="matrix(-1.4335232,0,0,1.4341698,269.48337,290.45712)" ns1:label="#g5607" id="default-pointer-c-1-2" style="display:inline">
        <ns0:path style="color:#000000;fill:url(#linearGradient4726-2-4-0);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.49009043;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 Z" id="path5565-2-4" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path ns2:nodetypes="cccccccc" id="path6242-4-9" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 Z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.49009043;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:0.98018089, 0.49009044;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:g transform="matrix(-1.4335232,0,0,1.4341698,311.05554,329.17971)" ns1:label="#g5607" id="default-pointer-c-1-2-5" style="display:inline">
        <ns0:path style="color:#000000;fill:url(#linearGradient4726-2-4-7-0);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.49009043;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 Z" id="path5565-2-4-9" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path ns2:nodetypes="cccccccc" id="path6242-4-9-7" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 Z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.49009043;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:0.98018089, 0.49009044;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g11020" transform="translate(-35,-4.36217)">
      <ns0:path transform="translate(2,453.36217)" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" ns2:ry="17" ns2:rx="17" ns2:cy="278" ns2:cx="120" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
      <ns0:text id="text11016" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan11018" ns2:role="line" style="font-size:14px;line-height:1.25">1</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g transform="translate(373,-4.36217)" id="g6104">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path6106" ns2:cx="120" ns2:cy="278" ns2:rx="17" ns2:ry="17" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" transform="translate(2,453.36217)"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" id="text6108"><ns0:tspan ns2:role="line" id="tspan6110" x="122.29289" y="736.36218" style="font-size:14px;line-height:1.25">2</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g id="g6112" transform="matrix(-1.4230531,0,0,1.4230531,989.7778,373.47398)">
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:2.10814333;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 146.93753,371.19797 0,-129.07529 143.35232,0" id="path6114" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
      <ns0:path id="path6116" style="fill:none;stroke:#000000;stroke-width:0.70271444px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" d="m 148.37105,270.089 c 0,-3.56432 2.88813,-6.45377 6.45085,-6.45377 l 156.25403,0" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
      <ns0:path id="path6122" style="fill:none;stroke:#000000;stroke-width:2.10814333;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 146.93753,270.089 c 0,-3.56432 2.88813,-6.45377 6.45085,-6.45377 l 82.9074,0" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
      <ns0:g style="display:inline" id="g6124" ns1:label="#g5607" transform="matrix(-1.4335232,0,0,1.4341698,-39.17119,345.97122)"/>
      <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1.06985807;marker:none;enable-background:accumulate" d="M 729.71875,115.75 718.1875,127.28125 H 571.125 c -5.55964,0 -10.03125,4.47161 -10.03125,10.03125 v 183.40625 c 0,5.55964 4.47161,10.0625 10.03125,10.0625 h 183.40625 c 5.55964,0 10.0625,-4.50286 10.0625,-10.0625 V 137.3125 c 0,-5.55964 -4.50286,-10.03125 -10.0625,-10.03125 h -13.3125 z" transform="matrix(-0.70271447,0,0,0.70271447,695.53118,187.29169)" id="rect6144" ns1:connector-curvature="0" ns2:nodetypes="ccsssssssscc"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:4.57940245;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect898" width="139.61769" height="21.314365" x="-299.73987" y="354.26465" transform="scale(-1,1)" rx="0" ry="0"/>
      <ns0:g ns1:label="pegged cogged wheel peg cog wood circle" id="g15931" style="display:inline;fill:#000000;enable-background:new" transform="matrix(-0.87496819,0,0,0.87496819,305.54804,-226.17153)">
        <ns0:title id="title15925">inställningar</ns0:title>
        <ns0:path ns1:connector-curvature="0" style="display:inline;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.06232423;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" d="m 367.48438,321.02344 c -0.55245,0 -0.99805,0.4456 -0.99805,0.99804 v 0.45118 a 5.7338295,5.73383 0 0 0 -1.35547,0.5664 l -0.32227,-0.32226 c -0.39063,-0.39064 -1.01952,-0.39064 -1.41015,0 l -0.70508,0.70508 c -0.39064,0.39062 -0.39064,1.01952 0,1.41015 l 0.32031,0.32031 a 5.7338295,5.73383 0 0 0 -0.56055,1.35743 H 362 c -0.55244,0 -0.99805,0.44365 -0.99805,0.99609 v 0.99805 c 0,0.55244 0.44561,0.99609 0.99805,0.99609 h 0.44922 a 5.7338295,5.73383 0 0 0 0.5664,1.35547 l -0.32226,0.32226 c -0.39064,0.39064 -0.39064,1.01953 0,1.41016 l 0.70508,0.70508 c 0.39063,0.39063 1.01952,0.39063 1.41015,0 l 0.32032,-0.32031 a 5.7338295,5.73383 0 0 0 1.35742,0.56054 v 0.45508 c 0,0.55244 0.4456,0.99609 0.99805,0.9961 h 0.99609 c 0.55244,0 0.99805,-0.44366 0.99805,-0.9961 v -0.45117 a 5.7338295,5.73383 0 0 0 1.35546,-0.56641 l 0.32227,0.32227 c 0.39064,0.39063 1.01952,0.39063 1.41016,0 l 0.70507,-0.70508 c 0.39064,-0.39063 0.39064,-1.01952 0,-1.41016 l -0.32031,-0.32031 A 5.7338295,5.73383 0 0 0 373.51172,329.5 h 0.45312 c 0.55245,0 0.99805,-0.44365 0.99805,-0.99609 v -0.99805 c 0,-0.55244 -0.4456,-0.99609 -0.99805,-0.99609 h -0.44922 a 5.7338295,5.73383 0 0 0 -0.5664,-1.35547 l 0.32226,-0.32227 c 0.39064,-0.39063 0.39064,-1.01953 0,-1.41015 l -0.70507,-0.70508 c -0.39064,-0.39064 -1.01952,-0.39064 -1.41016,0 l -0.32031,0.32031 a 5.7338295,5.73383 0 0 0 -1.35742,-0.56055 v -0.45508 c 0,-0.55244 -0.44561,-0.99804 -0.99805,-0.99804 z M 368,325 a 3,3 0 0 1 3,3 3,3 0 0 1 -3,3 3,3 0 0 1 -3,-3 3,3 0 0 1 3,-3 z" transform="translate(-348,348)" id="rect991-5"/>
      </ns0:g>
      <ns0:path ns1:connector-curvature="0" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1.40542889;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" d="m 265.54167,362.60228 v 23.57809 l -5.32168,-5.19732 -3.04096,6.21143 c -0.74485,1.67996 -4.61718,0.32918 -3.51611,-1.9173 l 3.00928,-6.44912 h -6.71545 z" id="path6128" ns2:nodetypes="cccccccc"/>
    </ns0:g>
    <ns0:g transform="translate(-388.97133,676.10528)" id="g12006">
      <ns0:g id="g5525" transform="translate(689,-168)" ns1:label="audio-volume-medium" style="display:inline">
        <ns0:path ns2:nodetypes="ccccccccc" id="path5533" d="m 20,222 2.484375,0 2.968754,-3 0.546871,0.0156 0,11 -0.475297,8.3e-4 L 22.484375,227 20,227 l 0,-5 z" style="color:#bebebe;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" ns1:connector-curvature="0"/>
        <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" id="rect5535" width="16" height="16" x="20" y="217" ns1:label="audio-volume-high"/>
        <ns0:path clip-path="url(#clipPath6279-7-9-7)" ns2:type="arc" style="fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path3718-5" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
        <ns0:path clip-path="url(#clipPath6265-3-4-4)" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3726-1" style="fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" ns2:type="arc" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
        <ns0:path clip-path="url(#clipPath6259-8-81-2)" ns2:type="arc" style="opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path3728-0" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
      </ns0:g>
      <ns0:g transform="translate(689,-639)" ns1:label="system-shutdown" id="g4692-3" style="display:inline">
        <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect10837-3-0" y="688" x="40" ry="0.15129246" rx="0.14408804" height="16" width="16"/>
        <ns0:path ns2:open="true" ns2:end="10.471045" ns2:start="5.239857" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" d="m 51.52343,689.95141 c 3.340544,1.94594 4.471097,6.23148 2.52516,9.57202 -1.945936,3.34054 -6.231476,4.4711 -9.57202,2.52516 -3.340544,-1.94594 -4.471097,-6.23148 -2.52516,-9.57202 0.612757,-1.05191 1.489249,-1.92583 2.542951,-2.53549" ns2:ry="7" ns2:rx="7" ns2:cy="696" ns2:cx="48" id="path3869-2" style="color:#000000;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
        <ns0:path ns2:nodetypes="cc" id="path4710" d="m 48,689 0,5" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:g id="g12661" transform="translate(666.07286,-166.91767)" ns1:label="network-wired" style="display:inline">
        <ns0:rect ns1:label="audio-volume-high" y="217" x="20" height="16" width="16" id="rect12673" style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible"/>
        <ns0:path id="rect12675" transform="translate(80,257)" d="m -55.25,-40 c -0.952203,0 -1.75,0.7978 -1.75,1.75 l 0,4.5 c 0,0.9522 0.797797,1.75 1.75,1.75 l 0.125,0 -0.78125,1.5625 -0.71875,1.4375 1.625,0 6,0 1.625,0 -0.71875,-1.4375 L -48.875,-32 l 0.125,0 c 0.952203,0 1.75,-0.7978 1.75,-1.75 l 0,-4.5 c 0,-0.9522 -0.797797,-1.75 -1.75,-1.75 l -6.5,0 z m 0.25,2 6,0 0,4 -6,0 0,-4 z" style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#bebebe;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans" ns1:connector-curvature="0"/>
        <ns0:path style="color:#bebebe;fill:none;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible" d="m 88,196 0,4" id="path12679" transform="translate(-60.0003,30)" ns1:connector-curvature="0"/>
        <ns0:path style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible" d="m 21.99975,231 12,0" id="path12681" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="rect12003" d="m 759.10724,57.4163 -3.74999,3.750004 -3.75001,-3.750005 z" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:g>
    <ns0:use x="0" y="0" ns4:href="#g12006" id="use15062" transform="translate(399,0)" width="840" height="400"/>
  </ns0:g>
</ns0:svg>
