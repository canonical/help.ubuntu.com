<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Klicka och flytta muspekaren med det numeriska tangentbordet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="a11y.html" title="Hjälpmedel">Hjälpmedel</a> › <a class="trail" href="a11y.html#mobility" title="Rörelsehinder">Rörelsehinder</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Klicka och flytta muspekaren med det numeriska tangentbordet</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du har svårt att använda en mus eller andra pekdon kan du styra musmarkören via det numeriska tangentbordet på ditt tangentbord. Denna funktion kallas <span class="em">mustangenter</span>.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps">
<p class="p">Öppna <span class="gui"><a href="shell-introduction.html#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Hjälpmedel</span>.</p>
<p class="p">Du kan nå översiktsvyn <span class="gui">Aktiviteter</span> genom att trycka på den, genom att flytta musmarkören till det övre, vänstra hörnet av skärmen, genom att trycka <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span> följt av <span class="key"><kbd>Retur</kbd></span> eller genom att trycka på <span class="key"><a href="keyboard-key-super.html" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span>.</p>
</li>
<li class="steps"><p class="p">Klicka på <span class="gui">Hjälpmedel</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Använd upp- och neråtpiltangenterna för att välja <span class="gui">Mustangenter</span> i avsnittet <span class="gui">Peka och klicka</span> och tryck sedan på <span class="key"><kbd>Retur</kbd></span> för att slå om <span class="gui">Mustangenter</span> till <span class="gui">På</span>.</p></li>
<li class="steps"><p class="p">Säkerställ att <span class="key"><kbd>Num Lock</kbd></span> är avstängd. Du kommer nu kunna flytta muspekaren med den numeriska delen av tangentbordet.</p></li>
</ol></div></div></div>
<p class="p">Det numeriska tangentbordet består av en mängd siffertangenter på ditt tangentbord, vanligtvis arrangerade som en fyrkant. Om du har ett tangentbord utan en numerisk del (som till exempel tangentbordet på en bärbar dator) kan du vara tvungen att hålla ner funktionstangenten (<span class="key"><kbd class="key-Fn">Fn</kbd></span>) och använda vissa andra knappar på ditt tangentbord som ett numeriskt tangentbord. Om du använder denna funktion ofta med en bärbar dator kan du köpa externa numeriska USB- eller Bluetooth-tangentbord.</p>
<p class="p">Varje siffra på det numeriska tangentbordet motsvarar en riktning. Till exempel om du trycker på <span class="key"><kbd>8</kbd></span> flyttar markören uppåt och om du trycker på <span class="key"><kbd>2</kbd></span> flyttar den neråt. Tryck på <span class="key"><kbd>5</kbd></span> för att klicka en gång med musen eller klicka på den två gånger snabbt för att dubbelklicka.</p>
<p class="p">De flesta tangentbord har en speciell tangent som låter dig högerklicka. Ibland kallas den <span class="key"><a href="keyboard-key-menu.html" title="Vad är Windows-tangenten?"><kbd>Meny</kbd></a></span>-tangenten. Notera dock att denna tangent reagerar på var tangentbordfokus är, inte var din musmarkör är. Se <span class="link"><a href="a11y-right-click.html" title="Simulera ett högerklick">Simulera ett högerklick</a></span> för information om hur du högerklickar genom att hålla ner <span class="key"><kbd>5</kbd></span> eller den vänstra musknappen.</p>
<p class="p">Om du vill använda det numeriska tangentbordet för att skriva siffror medan mustangenter är aktiverade, slå på <span class="key"><kbd>Num Lock</kbd></span>. Musen kan dock inte styras med det numeriska tangentbordet medan <span class="key"><kbd>Num Lock</kbd></span> är på.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">De normala siffertangenterna, i en rad i tangentbordets överkant, kommer inte styra muspekaren. Bara det numeriska tangentbordet kan användas till det här.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="mouse.html" title="Mus">Mus</a><span class="desc"> — <span class="link"><a href="mouse-lefthanded.html" title="Använd din mus med vänster hand">Vänsterhänt</a></span>, <span class="link"><a href="mouse-sensitivity.html" title="Justera hastigheten för musen och styrplattan">hastighet och känslighet</a></span>, <span class="link"><a href="mouse-touchpad-click.html" title="Klicka, dra eller rulla med styrplattan">klickning och rullning med styrplatta</a></span>…</span>
</li>
<li class="links "><a href="a11y.html#mobility" title="Rörelsehinder">Rörelsehinder</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
