<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skrivbord, program &amp; fönster</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Skrivbord, program &amp; fönster</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="whats-new.html" title="Vad är nytt i Ubuntu 14.04?"><span class="title">Vad är nytt i Ubuntu 14.04?</span><span class="linkdiv-dash"> — </span><span class="desc">Förbättringar i den senaste versionen av Ubuntu.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-introduction.html" title="Välkommen till Ubuntu"><span class="title">Välkommen till Ubuntu</span><span class="linkdiv-dash"> — </span><span class="desc">A visual introduction to the Unity desktop.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="shell-keyboard-shortcuts.html" title="Användbara kortkommandon"><span class="title">Användbara kortkommandon</span><span class="linkdiv-dash"> — </span><span class="desc">Get around the desktop using the keyboard.</span></a></div></div>
</div></div></div></div>
<div id="desktop" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Skrivbordet</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="unity-launcher-intro.html" title="Använda programstartaren"><span class="title">Använda programstartaren</span><span class="linkdiv-dash"> — </span><span class="desc">The Launcher is at the left of your screen.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen"><span class="title">Hantera program &amp; inställningar via menypanelen</span><span class="linkdiv-dash"> — </span><span class="desc">The menu bar is the dark strip on the top of your screen.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-dash-intro.html" title="Hitta program, filer, musik och annat med Dash"><span class="title">Hitta program, filer, musik och annat med Dash</span><span class="linkdiv-dash"> — </span><span class="desc">The Dash is the top button in the Launcher.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="clock-calendar.html" title="Kalendermöten"><span class="title">Kalendermöten</span><span class="linkdiv-dash"> — </span><span class="desc">Visa dina möten i kalendern överst i skärmen.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="unity-scrollbars-intro.html" title="What are overlay scrollbars?"><span class="title">What are overlay scrollbars?</span><span class="linkdiv-dash"> — </span><span class="desc">Overlay scrollbars are the thin orange strips on long documents.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-hud-intro.html" title="What is the HUD?"><span class="title">What is the HUD?</span><span class="linkdiv-dash"> — </span><span class="desc">Use the HUD to search menus of the apps you use.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-guest-session.html" title="Launch a restricted guest session"><span class="title">Launch a restricted guest session</span><span class="linkdiv-dash"> — </span><span class="desc">Let a friend or colleague borrow your computer in a secure manner.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-exit.html" title="Logga ut, stäng av, växla användare"><span class="title">Logga ut, stäng av, växla användare</span><span class="linkdiv-dash"> — </span><span class="desc">Learn how to leave your user account, by logging out, switching users,
    and so on.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="apps" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Program och fönster</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-apps-favorites.html" title="Change which applications show in the Launcher"><span class="title">Change which applications show in the Launcher</span><span class="linkdiv-dash"> — </span><span class="desc">Add, move, or remove frequently-used program icons on the 
    Launcher.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-windows.html" title="Fönster och arbetsytor"><span class="title">Fönster och arbetsytor</span><span class="linkdiv-dash"> — </span><span class="desc">Move and organize your windows.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="shell-windows-switching.html" title="Switch between windows"><span class="title">Switch between windows</span><span class="linkdiv-dash"> — </span><span class="desc">Press <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span>.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
