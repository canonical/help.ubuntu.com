<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>How do administrative privileges work?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="user-accounts.html" title="Användarkonton">Users</a> › <a class="trail" href="user-accounts.html#privileges" title="User privileges">Privileges</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">How do administrative privileges work?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">As well as the files that <span class="em">you</span> create, your computer has a number
 of files which are needed by the system for it to work properly. If these
 important <span class="em">system files</span> are changed improperly they can cause various
 things to break, so they are protected from changes by default. Certain
 applications also modify important parts of the system, and so are also
 protected.</p>
<p class="p">The way that they are protected is by only allowing users with
 <span class="em">administrative privileges</span> to change the files or use the applications.
 In day-to-day use, you won't need to change any system files or use these
 applications, so by default you do not have admin privileges.</p>
<p class="p">Sometimes you need to use these applications, so you may be able to
 temporarily get admin privileges to allow you to make the changes. If an
 application needs admin privileges, it will ask for your password. For example,
 if you want to install some new software, the software installer (package
 manager) will ask for your admin password so it can add the new application to
 the system. Once it has finished, your admin privileges will be taken away
 again.</p>
<p class="p">Admin privileges are associated with your user account. Some users are
 allowed to have admin privileges and some are not. Without admin privileges you
 will not be able to install software. Some user accounts (for example, the
 "root" account) have permanent admin privileges. You shouldn't use admin
 privileges all of the time, because you might accidentally change something
 you did not intend to (like delete a needed system file, for example).</p>
<p class="p">In summary, admin privileges allow you to change important parts of your
 system when needed, but prevent you from doing it accidentally.</p>
<div class="note" title="Anteckning"><div class="inner">
<div class="title title-note"><h2><span class="title">What does "super user" mean?</span></h2></div>
<div class="region"><div class="contents"><p class="p">A user with admin privileges is sometimes called a <span class="em">super user</span>.
 This is simply because that user has more privileges than normal users. You
 might see people discussing things like <span class="cmd">su</span> and <span class="cmd">sudo</span>;
 these are programs for temporarily giving you "super user" (admin) privileges.</p></div></div>
</div></div>
</div>
<div id="advantages" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Why are admin privileges useful?</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Requiring users to have admin privileges before important system changes
 are made is useful because it helps to prevent your system from being broken,
 intentionally or unintentionally.</p>
<p class="p">If you had admin privileges all of the time, you might accidentally change
 an important file, or run an application which changes something important by
 mistake. Only getting admin privileges temporarily, when you need them, reduces
 the risk of these mistakes happening.</p>
<p class="p">Only certain trusted users should be allowed to have admin privileges.
 This prevents other users from messing with the computer and doing things like
 uninstalling applications that you need, installing applications that you don't
 want, or changing important files. This is useful from a security standpoint.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="user-accounts.html#privileges" title="User privileges">User privileges</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="user-admin-change.html" title="Change who has administrative privileges">Change who has administrative privileges</a><span class="desc"> — You can change which users are allowed to make changes to the system
 by giving them administrative privileges.</span>
</li>
<li class="links ">
<a href="net-othersedit.html" title="Other users can't edit the network connections">Other users can't edit the network connections</a><span class="desc"> — You need to uncheck the <span class="gui">Available to all users</span> option in the network connection settings.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
