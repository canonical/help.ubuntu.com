<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Visuell överblick över GNOME</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 24.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Visuell överblick över GNOME</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">GNOME erbjuder ett användargränssnitt som designats för att inte vara i vägen, minimera distraktioner och hjälpa dig att få saker gjorda. När du loggar in första gången kommer du att se översiktsvyn <span class="gui">Aktiviteter</span> och systemraden.</p>
<div class="media media-image if-if if__not-target-mobile"><div class="inner"><img src="figures/shell-top-bar.png" width="600" class="media media-block" alt="GNOME-skalets systemrad"></div></div>
<p class="p">Systemraden erbjuder tillgång till dina fönster och program, din kalender och möten och <span class="link"><a href="status-icons.html.sv" title="Vad betyder ikonerna i systemraden?">systemegenskaper</a></span> som ljud, nätverk och ström. I systemmenyn i systemraden kan du ändra volym eller ljusstyrka för skärmen, redigera dina <span class="gui">Trådlösa</span> anslutningsdetaljer, kontrollera din batteristatus, logga ut eller växla användare och stänga av din dator.</p>
<div role="navigation" class="links sectionlinks"><div class="inner"><div class="region"><ul>
<li class="links "><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Översiktsvyn <span class="gui">Aktiviteter</span></a></li>
<li class="links "><a href="shell-introduction.html.sv#clock" title="Klocka, kalender och möten">Klocka, kalender och möten</a></li>
<li class="links "><a href="shell-introduction.html.sv#systemmenu" title="Systemmeny">Systemmeny</a></li>
<li class="links "><a href="shell-introduction.html.sv#lockscreen" title="Låsskärmen">Låsskärmen</a></li>
<li class="links "><a href="shell-introduction.html.sv#window-list" title="Fönsterlist">Fönsterlist</a></li>
</ul></div></div></div>
</div>
<section id="activities"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Översiktsvyn <span class="gui">Aktiviteter</span></span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Då du startar GNOME hamnar du automatiskt i översiktsvyn <span class="gui">Aktiviteter</span>. Översiktsvyn låter dig komma åt dina fönster och program. I översiktsvyn kan du också helt enkelt börja skriva för att söka bland dina program, filer, mappar och på webben.</p>
<p class="p">För att komma till översiktsvyn när som helst, klicka på knappen Aktiviteter i det övre vänstra hörnet eller flytta helt enkelt din muspekare till övre vänstra hörnet. Du kan också trycka på tangenten <span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span> på ditt tangentbord.</p>
<div class="media media-image floatend"><div class="inner"><img src="figures/shell-activities-dash.png" height="65" class="media media-block" alt="Activities button and Dash"></div></div>
<p class="p">Längst ner i översiktsvyn hittar du <span class="em">snabbstartspanelen</span>. Snabbstartspanelen visar dig dina favoritprogram och körande program. Klicka på vilken ikon som helst i favoriter för att öppna det programmet; om programmet redan körs kommer det att ha en liten punkt under sin ikon. Att klicka på dess ikon kommer att plocka fram det senast använda fönstret. Du kan också dra ikonen till en arbetsyta.</p>
<p class="p">Om du högerklickar på ikonen visas en meny som låter dig välja vilket fönster som helst för ett körande program, eller öppna ett nytt fönster. Du kan också klicka på ikonen medan du håller ner <span class="key"><kbd>Ctrl</kbd></span> för att öppna ett nytt fönster.</p>
<p class="p">När du går in i översiktsvyn kommer du först att hamna i fönsteröversiktsvyn. Denna visar dig live-uppdaterade miniatyrbilder av alla fönster på den aktuella arbetsytan.</p>
<p class="p">Klicka på rutnätsknappen (som har nio punkter) i snabbstartspanelen för att visa programöversiktsvyn. Denna visar dig alla program som finns installerade på din dator. Klicka på vilket program som helst för att köra det eller dra ett program till en arbetsyta som visas ovanför de installerade programmen. Du kan också dra ett program till snabbstartspanelen för att göra det till en favorit. Dina favoritprogram stannar kvar i snabbstartspanelen även om de inte kör, så att du kan nå dem snabbt.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="shell-apps-open.html.sv" title="Starta program">Läs mer om att starta program.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="shell-windows.html.sv" title="Fönster och arbetsytor">Läs mer om fönster och arbetsytor.</a></span></p></li>
</ul></div></div></div>
</div></div>
</div></section><section id="clock"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Klocka, kalender och möten</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="media media-image floatend if-if if__not-target-mobile"><div class="inner"><img src="figures/shell-appts.png" width="250" class="media media-block" alt="Klocka, kalender, möten och aviseringar"></div></div>
<p class="p">Klicka på klockan i systemraden för att se det aktuella datumet, en månadskalender och en lista på dina kommande möten och nya aviseringar. Du kan också öppna kalendern genom att trycka <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>V</kbd></span></span>. Du kan nå datum- och tidsinställningar och öppna hela ditt kalenderprogram direkt från menyn.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="clock-calendar.html.sv" title="Kalendermöten">Läs mer om kalendern och möten.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="shell-notifications.html.sv" title="Aviseringar och aviseringslistan">Läs mer om aviseringar och aviseringslistan.</a></span></p></li>
</ul></div></div></div>
</div></div>
</div></section><section id="systemmenu"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Systemmeny</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="media media-image floatend if-if if__not-target-mobile"><div class="inner"><img src="figures/shell-exit.png" width="250" class="media media-block" alt="Användarmeny"></div></div>
<p class="p">Klicka på systemmenyn i det övre högra hörnet för att hantera dina systeminställningar och din dator. Menyns övre del visar batteriets statusindikator och knappar för att starta Inställningar och skärmbildsverktyget. Knappen <span class="media"><span class="media media-image"><img src="figures/system-shutdown-symbolic.svg" class="media media-inline" alt="power"></span></span> låter dig försätta datorn i vänteläge eller slå av den, eller snabbt ge någon annan åtkomst till datorn utan att logga ut fullständigt. Skjutreglage låter dig styra systemvolymen eller skärmens ljusstyrka.</p>
<p class="p">Resten av menyn består av snabbinställningsknappar vilka låter dig snabbt styra tillgängliga tjänster och enheter såsom trådlöst nätverk, Bluetooth, ströminställningar och bakgrundsprogram.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="shell-exit.html.sv" title="Logga ut, stäng av eller växla användare">Läs mer om att växla användare, logga ut och stänga av din dator.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="quick-settings.html.sv" title="Snabbinställningar">Läs mer om snabbinställningar.</a></span></p></li>
</ul></div></div></div>
</div></div>
</div></section><section id="lockscreen"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Låsskärmen</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">När du låser din skärm eller den låses automatiskt så visas låsskärmen. Förutom att skydda ditt skrivbord medan du är borta från datorn så visar låsskärmen datum och tid. Den visar också information om din batteri- och nätverksstatus.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="shell-lockscreen.html.sv" title="Låsskärmen">Läs mer om låsskärmen.</a></span></p></li></ul></div></div></div>
</div></div>
</div></section><section id="window-list"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Fönsterlist</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">GNOME erbjuder ett annat sätt att växla mellan fönster än en permanent synlig fönsterlist som brukar finnas i andra skrivbordsmiljöer. Detta låter dig fokusera på dina uppgifter utan distraktioner.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="shell-windows-switching.html.sv" title="Växla mellan fönster">Läs mer om att växla fönster</a></span></p></li></ul></div></div></div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="shell-overview.html.sv" title="Ditt skrivbord">Ditt skrivbord</a><span class="desc"> — Arbeta med program, fönster och arbetsytor. Se dina möten och saker som är viktiga i systemraden.</span>
</li>
<li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
</ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
