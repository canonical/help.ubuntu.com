<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skriv speciella tecken</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="tips.html" title="Tips och tricks">Tips och tricks</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Skriv speciella tecken</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan skriva in och se tusentals tecken från de flesta av världens alla skrivsystem, även de som inte finns på ditt tangentbord. Den här sidan räknar upp några olika sätt för att skriva in specialtecken.</p>
<div role="navigation" class="links sectionlinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Metoder för att skriva in tecken</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="tips-specialchars.html#charmap" title="Teckenkarta">Teckenkarta</a></li>
<li class="links "><a href="tips-specialchars.html#ctrlshiftu" title="Kodpunkter">Kodpunkter</a></li>
<li class="links "><a href="tips-specialchars.html#sources" title="Inmatningskällor">Inmatningskällor</a></li>
</ul></div>
</div></div>
</div>
<div id="charmap" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Teckenkarta</span></h2></div>
<div class="region"><div class="contents">
<p class="p">GNOME inkluderar ett program med en teckenkarta som låter dig bläddra bland alla tecken i Unicode. Använd teckenkartan för att hitta tecknet du vill ha, och kopiera/klistra sedan in det där du vill ha det.</p>
<p class="p">Du kan hitta <span class="app">Teckenkarta</span> i <span class="gui">Snabbstartspanelen</span>. För mer information om teckenkartan, se <span class="link"><a href="https://help.gnome.org/users/gucharmap/stable/" title="https://help.gnome.org/users/gucharmap/stable/">handboken för Teckenkarta</a></span>.</p>
</div></div>
</div></div>
<div id="ctrlshiftu" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kodpunkter</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan skriva in Unicode-tecken med bara ditt tangentbord med tecknets numeriska kod. Varje tecken identifieras av en fyra tecken lång kod. För att hitta koden för ett tecken, hitta tecknet i teckenkartsprogrammet och titta i statusraden, eller i fliken <span class="gui">Teckendetaljer</span>. Koden är de fyra tecken som står efter <span class="gui">U+</span>.</p>
<p class="p">För att skriva in ett tecken med dess kod, tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>U</kbd></span></span>, skriv koden med fyra tecken, och tryck <span class="key"><kbd>Retur</kbd></span>. Om du ofta använder tecken som du inte enkelt kan komma åt med andra metoder kan du ha nytta av att memorera koden för dessa tecken så att du snabbt kan skriva in dem.</p>
</div></div>
</div></div>
<div id="sources" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Inmatningskällor</span></h2></div>
<div class="region"><div class="contents"><p class="p">Du kan ställa in att ditt tangentbord ska fungera som ett tangentbord för ett annat språk, oavsett vilka bokstäver som finns på tangenterna. Du kan också växla mellan olika inmatningskällor med en ikon i menyfältet. För att läsa mer, se <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">Använd alternativa inmatningskällor</a></span>.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="tips.html" title="Tips och tricks">Tips och tricks</a><span class="desc"> — <span class="link"><a href="tips-specialchars.html" title="Skriv speciella tecken">Speciella tecken</a></span>, <span class="link"><a href="mouse-middleclick.html" title="Mittenklick">mittenklick</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">Använd alternativa inmatningskällor</a><span class="desc"> — Lägg till indatakällor och växla mellan dem.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
