<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Filegenskaper</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Filegenskaper</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">För att visa information om en fil eller mapp, högerklicka på den och välj <span class="gui">Egenskaper</span>. Du kan också markera filen och trycka <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Retur</kbd></span></span>.</p>
<p class="p">Fönstret filegenskaper visa dig information som filtyp, filstorlek och när du senast modifierade den. Om du behöver denna information ofta kan du låta visa det i <span class="link"><a href="nautilus-list.html.sv" title="Kolumninställningar för listvy i Filer">listvykolumer</a></span> eller <span class="link"><a href="nautilus-display.html.sv#icon-captions" title="Ikonrubriker">ikonrubriker</a></span>.</p>
<p class="p">Informationen som finns på fliken <span class="gui">Grundläggande</span> förklaras nedan. De finns också flikar för <span class="gui"><span class="link"><a href="nautilus-file-properties-permissions.html.sv" title="Ange filrättigheter">Rättigheter</a></span></span> och <span class="gui"><span class="link"><a href="files-open.html.sv#default" title="Ändra standardprogrammet">Öppna med</a></span></span>. För vissa typer av filer, exempelvis för bilder och videor, så kommer det att finnas en extra flik med information så som dimensioner, längd och kodek.</p>
</div>
<div id="basic" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Grundläggande egenskaper</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Namn</span></dt>
<dd class="terms"><p class="p">Du kan byta namn på filen genom att ändra detta fält. Du kan också byta namn på en fil utanför egenskapsfönstret. Se <span class="link"><a href="files-rename.html.sv" title="Byt namn på en fil eller mapp">Byt namn på en fil eller mapp</a></span>.</p></dd>
<dt class="terms"><span class="gui">Typ</span></dt>
<dd class="terms">
<p class="p">Detta hjälper dig att identifiera filens typ, exempelvis PDF-dokument, OpenDocument-text eller JPEG-bild. Filtypen bestämmer bland annat vilket program som kan öppna filen. Du kan till exempel inte öppna en bild med en musikspelare. Se <span class="link"><a href="files-open.html.sv" title="Öppna filer med andra program">Öppna filer med andra program</a></span> för mer information om detta.</p>
<p class="p">Filens <span class="em">MIME-typ</span> visas i parenteser; MIME-typ är en standardmetod som datorer använder för att hänvisa till filtypen.</p>
</dd>
<dt class="terms">Innehåll</dt>
<dd class="terms"><p class="p">Det här fältet visas om du tittar på egenskaperna för en mapp istället för en fil. Det hjälper dig att se antal objekt i mappen. Om mappen innehåller andra mappar kommer varje underliggande mapp räknas som ett objekt, även om det innehåller andra objekt. Varje fil räknas också som ett objekt. Om mappen är tom kommer Innehåll visa <span class="gui">ingenting</span>.</p></dd>
<dt class="terms">Storlek</dt>
<dd class="terms">
<p class="p">Detta fält visas om du tittar på en fil (inte en mapp). Storleken för en fil berättar för dig hur mycket diskutrymme den upptar. Det är också en indikator på hur lång tid det tar att hämta ner en fil eller skicka den i ett e-postmeddelande (stora filer ta längre tid att skicka/ta emot).</p>
<p class="p">Storlekar kan anges i byte, KB, MB eller GB; i fallet med de sista tre så anges storleken i byte också inom parenteser. Tekniskt är 1KB 1024 byte, 1MB är 1024 KB och så vidare.</p>
</dd>
<dt class="terms">Föräldramapp</dt>
<dd class="terms"><p class="p">Platsen för varje fil på din dator anges av dess <span class="em">absoluta sökväg</span>. Detta är en unik ”adress” för filen på din dator, som utgörs av en lista av mappar som du måste gå in i för att hitta filen. Om Maria till exempel hade en fil som heter <span class="file">Resume.pdf</span> i sin Hemmapp, skulle dess föräldramapp bli <span class="file">/home/maria</span> och dess plats att bli <span class="file">/home/maria/Resume.pdf</span>.</p></dd>
<dt class="terms">Ledigt utrymme</dt>
<dd class="terms"><p class="p">Detta visas bara för mappar. Det visar hur mycket diskutrymme som finns tillgängligt på disken som mappen finns på. Detta gör det lättare att se om hårddisken är full.</p></dd>
<dt class="terms">Åtkommen</dt>
<dd class="terms"><p class="p">Tid och datum då filen senast öppnades.</p></dd>
<dt class="terms">Ändrad</dt>
<dd class="terms"><p class="p">Tid och datum när filen senast ändrades och sparades.</p></dd>
</dl></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html.sv#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="nautilus-file-properties-permissions.html.sv" title="Ange filrättigheter">Ange filrättigheter</a><span class="desc"> — Kontrollera vem som kan titta på och redigera dina filer och mappar.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
