<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Samba</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="version-control-ref.html" title="Referenser">Föregående</a><a class="nextlinks-next" href="samba-introduction.html" title="Inledning">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Samba</h1></div>
<div class="region">
<div class="contents"><p class="para">Datornätverk består ofta av flera olika system, och även om det vore trevligt att administrera ett nätverk som endast bestod av skrivbordsdatorer och servrar med Ubuntu måste somliga nätverk bestå av både Ubuntusystem och <span class="trademark">Microsoft®</span><span class="trademark">Windows®</span>-system som arbetar tillsammans i harmoni. Den här sektionen av <span class="phrase">Ubuntus</span> serverguide introducerar principer och verktyg som används till att konfigurera din Ubuntuserver till att dela nätverksresurser med Windowsdatorer.</p></div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="samba-introduction.html" title="Inledning">Inledning</a></li>
<li class="links"><a class="xref" href="samba-fileserver.html" title="File Server">File Server</a></li>
<li class="links"><a class="xref" href="samba-printserver.html" title="Skrivarserver">Skrivarserver</a></li>
<li class="links"><a class="xref" href="samba-fileprint-security.html" title="Securing File and Print Server">Securing File and Print Server</a></li>
<li class="links"><a class="xref" href="samba-dc.html" title="As a Domain Controller">As a Domain Controller</a></li>
<li class="links"><a class="xref" href="samba-ad-integration.html" title="Active Directory Integration">Active Directory Integration</a></li>
</ul></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="version-control-ref.html" title="Referenser">Föregående</a><a class="nextlinks-next" href="samba-introduction.html" title="Inledning">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
