<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Dölj en fil</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#faq" title="Tips och frågor">Tips och frågor</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Dölj en fil</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">GNOMEs filhanterare gör dig möjligheten att dölja och visa filer med ett enkelt kommando. När en fil är dold syns den inte i filhanteraren, men finns fortfarande i mappen.</p>
<p class="p">För att dölja en fil, <span class="link"><a href="files-rename.html" title="Byt namn på en fil eller mapp">döp om den</a></span> med en <span class="key"><kbd>.</kbd></span> i början av filnamnet. Exempel: För att dölja en fil med namnet <span class="file">exempel.txt</span> kan du döpa om den till <span class="file">.exempel.txt</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan dölja mappar på samma sätt som du döljer filer. Dölj en mapp genom att placera en <span class="key"><kbd>.</kbd></span> i början av mappens namn.</p></div></div></div></div>
</div>
<div id="show-hidden" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Visa alla dolda filer</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Om du vill se alla dolda filer i en mapp, gå till den mappen och klicka antingen på <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="nerknappen"></span></span> i verktygsraden och välj <span class="gui">Visa dolda filer</span> eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>H</kbd></span></span>. Du kommer se alla dolda filer, tillsammans med vanliga filer som inte är dolda.</p>
<p class="p">För att dölja filerna igen, klicka antingen på <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="nerknappen"></span></span> i verktygsraden och välj (avbocka) <span class="gui">Visa dolda filer</span> eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>H</kbd></span></span> igen.</p>
</div></div>
</div></div>
<div id="unhide" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Sluta dölja en fil</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att sluta dölja en fil, gå till mappen där filen finns och klicka på <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="nerknappen"></span></span> i verktygsraden och välj <span class="gui">Visa dolda filer</span>. Leta sedan upp den dolda filen och döp om den så att den inte har en <span class="key"><kbd>.</kbd></span> framför sitt namn. Exempel: För att sluta dölja en fil som heter <span class="file">.exempel.txt</span> bör du döpa om den till <span class="file">exempel.txt</span>.</p>
<p class="p">När du har döpt om filen kan du antingen klicka på <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="nerknappen"></span></span> i verktygsraden och välj <span class="gui">Visa dolda filer</span>, eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>H</kbd></span></span> för att dölja de andra dolda filerna igen.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Som standard ser du bara dolda filer i filhanteraren tills du stänger filhanteraren. För att ändra den inställningen så att filhanteraren alltid visar dolda filer, se <span class="link"><a href="nautilus-views.html" title="Visningsinställningar i Filer">Visningsinställningar i <span class="app">Filer</span></a></span>.</p></div></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">De flesta dolda filer har en <span class="key"><kbd>.</kbd></span> i början av filnamnet, men andra kan ha en <span class="key"><kbd>~</kbd></span> i slutet av filnamnet istället. Dessa filer är säkerhetskopior. Se <span class="link"><a href="files-tilde.html" title='Vad är en fil med ett "~" i slutet av filnamnet?'>Vad är en fil med ett "~" i slutet av filnamnet?</a></span> för mer information.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html#faq" title="Tips och frågor">Tips och frågor</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-tilde.html" title='Vad är en fil med ett "~" i slutet av filnamnet?'>Vad är en fil med ett "~" i slutet av filnamnet?</a><span class="desc"> — Detta är säkerhetskopior. De är dolda som standard.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
