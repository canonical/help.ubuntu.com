<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>What are overlay scrollbars?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Desktop</a> › <a class="trail" href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">What are overlay scrollbars?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Ubuntu includes <span class="em">overlay scrollbars</span> which take up less screen space than
traditional scrollbars, giving you more room for your content. While inspired by mobile devices
where traditional scrollbars aren't needed, Ubuntu's overlay scrollbars are designed to work
just as well with a mouse.</p>
<p class="p">Some apps like Firefox and LibreOffice don't support the new scrollbars yet.</p>
</div>
<div id="using" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Use the scrollbars</span></h2></div>
<div class="region"><div class="contents">
<p class="p">The overlay scrollbar appears as a thin orange strip at the edge of a scrollable area.
  The position of the scrollbar corresponds with your screen's position in the scrollable content.
  The strip length corresponds with the content length; the shorter the strip, the longer the content.</p>
<p class="p">Move your mouse pointer over any point on the scrollable edge of the content to reveal the <span class="gui">thumb slider</span>.</p>
<div class="list"><div class="inner">
<div class="title title-list"><h3><span class="title">Ways to use the scrollbars:</span></h3></div>
<div class="region"><ul class="list">
<li class="list"><p class="p">
    Click the top half of the <span class="gui">thumb slider</span> to scroll one page up. Click the bottom half to scroll one page down.
    </p></li>
<li class="list"><p class="p">
    Drag the <span class="gui">thumb slider</span> up or down to move the screen's position exactly where you want it.
    </p></li>
<li class="list"><p class="p">
    <span class="link"><a href="mouse-middleclick.html" title="Mittenklick">Mittenklick</a></span> on the <span class="gui">thumb slider</span> to move the screen's position without needing to drag or
    scroll page by page. This is especially useful in long documents.
    </p></li>
</ul></div>
</div></div>
</div></div>
</div></div>
<div id="disable-scrollbars" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Disable the scrollbars</span></h2></div>
<div class="region"><div class="contents">
<p class="p">You can disable the new scrollbars if you prefer the traditional style:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Open the <span class="app">Terminal</span> by pressing <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>t</kbd></span></span>
    or by searching for <span class="input">terminal</span> in the <span class="gui">Dash</span>.
    </p></li>
<li class="steps">
<p class="p">Type the following command and press <span class="key"><kbd>Enter</kbd></span>:</p>
<div class="code"><pre class="contents ">gsettings set com.canonical.desktop.interface scrollbar-mode normal</pre></div>
</li>
</ol></div></div></div>
<p class="p">If you change your mind and want to re-enable the scrollbars, run this command:</p>
<div class="code"><pre class="contents ">gsettings reset com.canonical.desktop.interface scrollbar-mode</pre></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Setting your theme to <span class="link"><a href="a11y-contrast.html" title="Justera kontrasten">High Contrast</a></span> will also disable the overlay scrollbars.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="mouse-touchpad-click.html" title="Klicka, dra, eller rulla med styrplattan">Klicka, dra, eller rulla med styrplattan</a><span class="desc"> — Klicka, dra, eller rulla genom att peta och använda gester på din styrplatta.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
