<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Why won't my computer turn back on after I suspended it?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="power.html#problems" title="Problem">Power problems</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="hardware-problems-graphics.html" title="Skärmproblem">Skärmproblem</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Why won't my computer turn back on after I suspended it?</span></h1></div>
<div class="region">
<div class="contents"><p class="p">If you <span class="link"><a href="power-suspend.html" title="What happens when I suspend my computer?">suspend</a></span> or <span class="link"><a href="power-hibernate.html" title="How do I hibernate my computer?">hibernate</a></span> your computer, then try to resume it or
turn it back on, you may find that it does not work as you expected. This could
be because suspend and hibernate aren't supported properly by your
hardware.</p></div>
<div id="resume" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">My computer is suspended and isn't resuming</span></h2></div>
<div class="region"><div class="contents">
<p class="p">If you suspend your computer and then press a key or click the mouse, it
  should wake up and display a screen asking for your password. If this doesn't
 happen, try pressing the power button (don't hold it in, just press it
  once).</p>
<p class="p">If this still doesn't help, make sure that your computer's monitor is
  switched on and try pressing a key on the keyboard again.</p>
<p class="p">As a last resort, turn off the computer by holding in the power button for
  5-10 seconds, although you will lose any unsaved work by doing this. You
  should then be able to turn on the computer again.</p>
<p class="p">If this happens every time you suspend your computer, the suspend
  feature may not work with your hardware.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">If your computer loses power and doesn't have an alternative power
    supply (such as a working battery), it will switch off.</p></div></div></div></div>
</div></div>
</div></div>
<div id="hibernate" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">None of my applications/documents are open when I turn on the computer
  again</span></h2></div>
<div class="region"><div class="contents">
<p class="p">If you hibernated your computer and switched it on again, but none of your
  documents or applications are open, it probably failed to hibernate properly.
  Sometimes this happens because of a minor problem, and the computer will be
  able to hibernate properly the next time you do it. It might also happen
  because you had installed a software update which required the computer to be
  restarted; in this case, the computer may have shut down instead of
  hibernating.</p>
<p class="p">It is also possible that the computer is not capable of hibernating
  because the hardware doesn't support it properly. This might be because of a
  problem with Linux drivers for your hardware, for example. You can test this
  by hibernating again and seeing if it works the second time. If it doesn't,
  it is probably a problem with your computer's drivers.</p>
</div></div>
</div></div>
<div id="hardware" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">My wireless connection (or other hardware) doesn't work when I wake
  up my computer</span></h2></div>
<div class="region"><div class="contents">
<p class="p">If you suspend or hibernate your computer and then resume it again, you
  may find that your internet connection, mouse, or some other device doesn't
  work properly. This could be because the device's driver doesn't
  properly support suspend or hibernate. This is a <span class="link"><a href="hardware-driver.html" title="Vad är en drivrutin?">problem with the driver</a></span> and not the device
  itself.</p>
<p class="p">If the device has a power switch, try turning it off and then on again. In
  most cases, the device will start working again. If it connects via a USB
  cable or similar, unplug the device and then plug it in again and see if it
  works.</p>
<p class="p">If you cannot turn off/unplug the device, or if this does not work, you
  may need to restart your computer for the device to start working again.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="power.html#problems" title="Problem">Power problems</a><span class="desc"> — Troubleshoot problems with power and batteries.</span>
</li>
<li class="links ">
<a href="hardware-problems-graphics.html" title="Skärmproblem">Skärmproblem</a><span class="desc"> — Felsök skärm- och grafikproblem.</span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="power-hibernate.html" title="How do I hibernate my computer?">How do I hibernate my computer?</a><span class="desc"> — Hibernate is disabled by default since it's not well supported.</span>
</li>
<li class="links ">
<a href="power-nowireless.html" title="I have no wireless network when I wake up my computer">I have no wireless network when I wake up my computer</a><span class="desc"> — Some wireless devices have problems handling when your computer is suspended and doesn't resume properly.</span>
</li>
<li class="links ">
<a href="power-closelid.html" title="Why does my computer turn off when I close the lid?">Why does my computer turn off when I close the lid?</a><span class="desc"> — Laptops go to sleep when you close the lid, in order to save power.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
