<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Staying safe on the internet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-general.html" title="Networking terms &amp; tips">Networking terms &amp; tips</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Staying safe on the internet</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">A possible reason for why you are using Ubuntu is the robust security that Linux based
systems are known for. One reason that Linux is relatively safe from malware and
viruses is due to the lower number of people who use it.
Viruses are targeted at popular operating systems like Windows, that have an extremely large
user base. Linux based systems are also very secure due to their open source nature, which allows
experts to modify and enhance the security features included with each distribution.</p>
<p class="p">Despite the measures taken to ensure that your installation of Ubuntu is secure, there
are always vulnerabilities. As an average user on the internet you can still be susceptible to:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Phishing Scams (websites and emails that try to obtain sensitive information through deception)</p></li>
<li class="list"><p class="p"><span class="link"><a href="net-email-virus.html" title="Do I need to scan my emails for viruses?">Forwarding malicious emails</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="net-antivirus.html" title="Behöver jag ett anti-virusprogram?">Applications with malicious intent (viruses)</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?">Unauthorized remote/local network access</a></span></p></li>
</ul></div></div></div>
<p class="p">To stay safe online, keep in mind the following tips:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Be wary of emails, attachments, or links that were sent from people you do not know.</p></li>
<li class="list"><p class="p">If a website's offer is too good to be true, or asks for sensitive information
that seems unnecessary, then think twice about what information you are submitting and the potential
consequences if that information is compromised by identity thieves or other criminals.</p></li>
<li class="list"><p class="p">Be careful in providing any application <span class="link"><a href="user-admin-explain.html" title="How do administrative privileges work?">root level permissions</a></span>, especially ones that
you have not used before or apps that are not well-known. Providing anyone/anything with root level
permissions puts your computer at high risk to exploitation.</p></li>
<li class="list"><p class="p">Make sure you are only running necessary remote-access services. Having
SSH or VNC running can be useful, but also leaves your computer open to intrusion if not
secured properly. Consider using a <span class="link"><a href="net-firewall-on-off.html" title="Enable or block firewall access">firewall</a></span> to help
protect your computer from intrusion.</p></li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-general.html" title="Networking terms &amp; tips">Networking terms &amp; tips</a><span class="desc"> — 
      <span class="link"><a href="net-findip.html" title="Hitta din IP-adress">Find your IP address</a></span>,
      <span class="link"><a href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?">WEP &amp; WPA security</a></span>,
      <span class="link"><a href="net-macaddress.html" title="What is a MAC address?">MAC addresses</a></span>,
      <span class="link"><a href="net-proxy.html" title="Define proxy settings">proxies</a></span>…
    </span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
