<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Trådlösa nätverk</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="net.html" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Trådlösa nätverk</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="net-wireless-connect.html" title="Anslut till ett trådlöst nätverk"><span class="title">Anslut till ett trådlöst nätverk</span><span class="linkdiv-dash"> — </span><span class="desc">Nå internet - trådlöst.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-manual.html" title="Ange nätverksinställningar manuellt"><span class="title">Ange nätverksinställningar manuellt</span><span class="linkdiv-dash"> — </span><span class="desc">Du kan behöva mata in nätverksinställningar om de inte tilldelas automatiskt.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-vpn-connect.html" title="Anslut till ett VPN"><span class="title">Anslut till ett VPN</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in en VPN-anslutning till ett lokalt nätverk över internet.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-hidden.html" title="Anslut till ett dolt, trådlöst nätverk"><span class="title">Anslut till ett dolt, trådlöst nätverk</span><span class="linkdiv-dash"> — </span><span class="desc">Anslut till ett trådlöst nätverk som inte visas i nätverkslistan.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-mobile.html" title="Anslut till mobilt bredband"><span class="title">Anslut till mobilt bredband</span><span class="linkdiv-dash"> — </span><span class="desc">Använd din telefon- eller internet-sticka för att ansluta till mobilt bredbandsnätverk.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-troubleshooting.html" title="Felsökning av trådlösa nätverk"><span class="title">Felsökning av trådlösa nätverk</span><span class="linkdiv-dash"> — </span><span class="desc">Identifiera och fixa problem med trådlösa anslutningar.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="net-wireless-noconnection.html" title="Jag har matat in rätt lösenord, men kan fortfarande inte ansluta"><span class="title">Jag har matat in rätt lösenord, men kan fortfarande inte ansluta</span><span class="linkdiv-dash"> — </span><span class="desc">Dubbelkolla lösenordet och andra saker att prova.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-find.html" title="Jag kan inte se mitt trådlösa nätverk i listan"><span class="title">Jag kan inte se mitt trådlösa nätverk i listan</span><span class="linkdiv-dash"> — </span><span class="desc">Det trådlösa nätverket kan vara avstängt eller trasigt eller så kan du försöka ansluta till ett dolt nätverk.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-adhoc.html" title="Skapa en trådlös surfzon"><span class="title">Skapa en trådlös surfzon</span><span class="linkdiv-dash"> — </span><span class="desc">Använd ett ad-hoc-nätverk för att låta andra enheter ansluta till din dator och dess nätverksanslutningar.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-airplane.html" title="Stäng av trådlöst (flygplansläge)"><span class="title">Stäng av trådlöst (flygplansläge)</span><span class="linkdiv-dash"> — </span><span class="desc">Öppna nätverksinställningar och slå om flygplansläge till PÅ.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-wepwpa.html" title="Vad betyder WEP och WPA?"><span class="title">Vad betyder WEP och WPA?</span><span class="linkdiv-dash"> — </span><span class="desc">WEP och WPA är sätt att kryptera data på trådlösa nätverk.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-disconnecting.html" title="Varför kopplar mitt trådlösa nätverk ner hela tiden?"><span class="title">Varför kopplar mitt trådlösa nätverk ner hela tiden?</span><span class="linkdiv-dash"> — </span><span class="desc">Du kan ha låg signal eller så kanske nätverket inte låter dig ansluta ordentligt.</span></a></div>
</div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a><span class="desc"> — <span class="link"><a href="net-wireless.html" title="Trådlösa nätverk">Trådlöst</a></span>, <span class="link"><a href="net-wired.html" title="Trådbundna nätverk">trådbundet</a></span>, <span class="link"><a href="net-problem.html" title="Nätverksproblem">anslutningsproblem</a></span>, <span class="link"><a href="net-browser.html" title="Webbläsare">webbsurfning</a></span>, <span class="link"><a href="net-email.html" title="E-post &amp; e-postprogramvara">e-postkonton</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="net-problem.html" title="Nätverksproblem">Nätverksproblem</a><span class="desc"> — <span class="link"><a href="net-wireless-troubleshooting.html" title="Felsökning av trådlösa nätverk">Felsök trådlösa anslutningar</a></span>, <span class="link"><a href="net-wireless-find.html" title="Jag kan inte se mitt trådlösa nätverk i listan">hitta ditt trådlösa nätverk</a></span>…</span>
</li>
<li class="links ">
<a href="net-general.html" title="Nätverkstermer &amp; -tips">Nätverkstermer &amp; -tips</a><span class="desc"> — <span class="link"><a href="net-findip.html" title="Hitta din IP-adress">Hitta din IP-adress</a></span>, <span class="link"><a href="net-wireless-wepwpa.html" title="Vad betyder WEP och WPA?">WEP- &amp; WPA-säkerhet</a></span>, <span class="link"><a href="net-macaddress.html" title="Vad är en MAC-adress?">MAC-adresser</a></span>, <span class="link"><a href="net-proxy.html" title="Definiera proxyinställningar">proxyservrar</a></span>…</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
