<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Kopiera eller flytta filer och mappar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#common-file-tasks" title="Vanliga åtgärder">Vanliga åtgärder</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Kopiera eller flytta filer och mappar</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">En fil eller mapp kan kopieras eller flyttas till en ny plats genom att dra och släppa den med musen, använda kommandona kopiera och klistra in eller via snabbtangenter.</p>
<p class="p">Du kanske vill kopiera en presentation till en minnessticka så du kan ta arbetet med dig. Eller så kan du göra en säkerhetskopia av ett dokument innan du gör ändringar i det (och sedan använda den gamla kopia om du inte tyckte om ändringarna).</p>
<p class="p">Dessa instruktioner gäller både filer och mappar. Du kopierar och flyttar filer och mappar på exakt samma sätt.</p>
<div class="steps ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-steps"><h2><span class="title">Kopiera och klistra in filer</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Markera den fil du vill kopiera genom att klicka på den en gång.</p></li>
<li class="steps"><p class="p">Högerklicka och välj <span class="gui">Kopiera</span>, eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>C</kbd></span></span>.</p></li>
<li class="steps"><p class="p">Navigera till en annan mapp, där du vill lägga kopian av filen.</p></li>
<li class="steps"><p class="p">Klicka på menyknappen och välj <span class="gui">Klistra in</span> för att kopiera filen, eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>V</kbd></span></span>. Det kommer nu att finnas en kopia av filen i originalmappen och den andra mappen.</p></li>
</ol></div>
</div>
</div>
<div class="steps ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-steps"><h2><span class="title">Klipp ut och klistra in filer för att flytta dem</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Markera filen du vill flytta genom att klicka på den en gång.</p></li>
<li class="steps"><p class="p">Högerklicka och välj <span class="gui">Klipp ut</span>, eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>X</kbd></span></span>.</p></li>
<li class="steps"><p class="p">Navigera till den mapp dit du vill flytta filen.</p></li>
<li class="steps"><p class="p">Klicka på menyknappen i verktygsfältet och välj <span class="gui">Klistra in</span> för att flytta filen, eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>V</kbd></span></span>. Filen kommer att tas från sin originalmapp och flyttas till den andra mappen.</p></li>
</ol></div>
</div>
</div>
<div class="steps ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-steps"><h2><span class="title">Dra filer för att kopiera eller flytta</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna filhanteraren och gå till mappen som innehåller filen du vill kopiera.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Filer</span> i systemraden och välj <span class="gui">Nytt fönster</span> (eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>N</kbd></span></span>) för att öppna ett andra fönster. I det nya fönstret, navigera till mappen där du önskar att flytta eller kopiera filen.</p></li>
<li class="steps">
<p class="p">Klicka och dra filen från ett fönster till det andra. Detta kommer att <span class="em">flytta den</span> om destinationen är på <span class="em">samma</span> enhet, eller <span class="em">kopiera den</span> om destinationen är på en <span class="em">annan</span> enhet.</p>
<p class="p">Om du till exempel drar en fil från en USB-minne till din Hemmapp kommer den att kopieras eftersom du drar den från en enhet till en annan.</p>
<p class="p">Du kan tvinga filen att kopieras genom att hålla ner tangenten <span class="key"><kbd>Ctrl</kbd></span> medan du drar eller tvinga den att flyttas genom att hålla ner tangenten <span class="key"><kbd>Skift</kbd></span> medan du drar.</p>
</li>
</ol></div>
</div>
</div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan inte kopiera eller flytta en fil in i en mapp som är <span class="em">skrivskyddad</span>. Vissa mappar är skrivskyddade för att förhindra att du gör ändringar i deras innehåll. Du kan ändra saker från att vara skrivskyddade genom att <span class="link"><a href="nautilus-file-properties-permissions.html.sv" title="Ange filrättigheter">ändra filrättigheterna</a></span>.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html.sv#common-file-tasks" title="Vanliga åtgärder">Vanliga åtgärder</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-browse.html.sv" title="Bläddra bland filer och mappar">Bläddra bland filer och mappar</a><span class="desc"> — Hantera och organisera filer med filhanteraren.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
