<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Handbok för Ubuntu-skrivbordet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" class="media media-inline" alt="Ubuntu Logo"></span></span> Handbok för Ubuntu-skrivbordet</span></h1></div>
<div class="region"><div class="contents">
<div class="links topiclinks"><div class="inner"><div class="region">
<div class="mouseovers"><img src="figures/unity.png"></div>
<ul class="mouseovers">
<li class="links"><a class="bold" href="whats-new.html" title="Vad är nytt i Ubuntu 14.04?">Vad är nytt i Ubuntu 14.04?</a></li>
<li class="links"><a class="bold" href="unity-introduction.html" title="Välkommen till Ubuntu"><img src="figures/ubuntu-mascot-creature.jpg">Välkommen till Ubuntu</a></li>
<li class="links"><a class="bold" href="unity-launcher-intro.html" title="Använda programstartaren"><img src="figures/unity-launcher-intro.png">Använda programstartaren</a></li>
<li class="links"><a class="bold" href="unity-dash-intro.html" title="Hitta program, filer, musik och annat med Dash"><img src="figures/unity-dash-intro.png">Hitta program, filer, musik och annat med Dash</a></li>
<li class="links"><a class="bold" href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen"><img src="figures/unity-appmenu-intro.png">Hantera program &amp; inställningar via menypanelen</a></li>
<li class="links"><a class="bold" href="shell-exit.html" title="Logga ut, stäng av, växla användare"><img src="figures/unity-exit.png">Logga ut, stäng av, växla användare</a></li>
</ul>
<div class="clear"></div>
</div></div></div>
<div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-grid ">
<div class="links-grid-link"><a href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord, program &amp; fönster</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="unity-introduction.html" title="Välkommen till Ubuntu">Introduktion</a></span>, <span class="link"><a href="shell-keyboard-shortcuts.html" title="Användbara kortkommandon">kortkommandon</a></span>, <span class="link"><a href="shell-windows.html" title="Fönster och arbetsytor">fönster</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="net-wireless.html" title="Trådlös anslutning">Trådlöst</a></span>, <span class="link"><a href="net-wired.html" title="Trådbunden anslutning">trådbundet</a></span>, <span class="link"><a href="net-problem.html" title="Nätverksproblem">anslutnings-problem</a></span>, <span class="link"><a href="net-browser.html" title="Webbläsare">webbnavigering</a></span>, <span class="link"><a href="net-email.html" title="E-post &amp; e-postmjukvara">e-postkonton</a></span>, <span class="link"><a href="net-chat.html" title="Chatt &amp; sociala medier">snabbmeddelanden</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="media.html#photos" title="Foton och digitalkameror">Digitala kameror</a></span>, <span class="link"><a href="media.html#music" title="Musik och bärbara ljudspelare">iPod-spelare</a></span>, <span class="link"><a href="media.html#videos" title="Videor och videokameror">spela upp videofilmer</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="addremove.html" title="Lägg till &amp; ta bort mjukvara">Lägg till &amp; ta bort mjukvara</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="addremove-install.html" title="Installera fler program">Installera</a></span>, <span class="link"><a href="addremove-remove.html" title="Ta bort ett program">ta bort</a></span>, <span class="link"><a href="addremove-sources.html" title="Lägg till fler programförråd">extra förråd</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="prefs.html" title="Inställningar för användare och system">Inställningar för användare och system</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html" title="Användarkonton">användarkonton</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="hardware.html" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="hardware.html#problems" title="Vanliga problem">Hårdvaruproblem</a></span>, <span class="link"><a href="printing.html" title="Utskrifter">skrivare</a></span>, <span class="link"><a href="power.html" title="På/av &amp; batteri">på/av-funktioner</a></span>, <span class="link"><a href="color.html" title="Hantera färginställningar">färginställningar</a></span>, <span class="link"><a href="bluetooth.html" title="Bluetooth">Bluetooth</a></span>, <span class="link"><a href="disk.html" title="Hårddiskar &amp; lagring">hårddiskar</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="a11y.html" title="Hjälpmedel">Hjälpmedel</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="a11y.html#vision" title="Synnedsättning">Syn</a></span>, <span class="link"><a href="a11y.html#sound" title="Hörselnedsättning">hörsel</a></span>, <span class="link"><a href="a11y.html#mobility" title="Rörelsehinder">rörlighet</a></span>, <span class="link"><a href="a11y-braille.html" title="Läs skärmen med punktskrift">punktskrift</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="tips.html" title="Tips och tricks">Tips och tricks</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="tips-specialchars.html" title="Skriv speciella tecken">Speciella tecken</a></span>, <span class="link"><a href="mouse-middleclick.html" title="Mittenklick">mittenklick</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="more-help.html" title="Få mer hjälp">Få mer hjälp</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="about-this-guide.html" title="Om denna handbok">Användningstips</a></span>, <span class="link"><a href="get-involved.html" title="Medverka till att förbättra den här handboken">hjälp till att förbättra handboken</a></span>…</span></div>
</div>
</div></div></div>
</div></div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
