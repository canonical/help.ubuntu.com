<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Jag kan inte ansluta min Bluetooth-enhet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html.sv#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="bluetooth.html.sv#problems" title="Problem">Bluetooth-problem</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Jag kan inte ansluta min Bluetooth-enhet</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Det finns ett flertal anledningar till varför du kanske inte kan ansluta till en Bluetooth-enhet, så som en telefon eller en hörlur.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Anslutning blockerad eller otillförlitlig</dt>
<dd class="terms"><p class="p">Vissa Bluetooth-enheter blockerar anslutningar som standard eller kräver att du ändrar en inställning för att tillåta anslutningar. Försäkra att din enhet är inställd för att tillåta anslutningar.</p></dd>
<dt class="terms">Bluetooth-hårdvara kändes inte igen</dt>
<dd class="terms"><p class="p">Din Bluetooth-adapter kanske inte har känts igen av datorn. Detta skulle kunna vara för att <span class="link"><a href="hardware-driver.html.sv" title="Vad är en drivrutin?">drivrutiner</a></span> för adaptern inte installerats. Vissa Bluetooth-adaptrar saknar stöd under Linux, så du kan kanske inte få tag i rätt drivrutiner för dessa. Om det är fallet kommer du troligtvis att behöva skaffa en annan Bluetooth-adapter.</p></dd>
<dt class="terms">Adaptern är inte påslagen</dt>
<dd class="terms"><p class="p">Försäkra att din Bluetooth-adapter är påslagen. Öppna Bluetooth-panelen och kontrollera att den inte är <span class="link"><a href="bluetooth-turn-on-off.html.sv" title="Aktivera eller inaktivera Bluetooth">inaktiverad</a></span>.</p></dd>
<dt class="terms">Enhetens Bluetooth-anslutning är avslagen</dt>
<dd class="terms"><p class="p">Kontrollera att Bluetooth är påslaget i enheten du försöker ansluta till och att den är <span class="link"><a href="bluetooth-visibility.html.sv" title="Vad är Bluetooth-synlighet?">detekterbar eller synlig</a></span>. Om du till exempel försöker ansluta till en telefon, säkerställ att den inte är i flygplansläge.</p></dd>
<dt class="terms">Ingen Bluetooth-adapter i din dator</dt>
<dd class="terms"><p class="p">Många datorer har inte Bluetooth-adaptrar. Du kan köpa en adapter om du vill använda Bluetooth.</p></dd>
</dl></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="bluetooth.html.sv#problems" title="Problem">Bluetooth-problem</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="hardware-driver.html.sv" title="Vad är en drivrutin?">Vad är en drivrutin?</a><span class="desc"> — En hårdvaru-/enhetsdrivrutin låter din dator använda enheter som ansluts till den.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p>You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
