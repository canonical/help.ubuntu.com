<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Time Synchronisation</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="networking.html" title="Nätverk">Nätverk</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="dhcp.html" title="Dynamic Host Configuration Protocol (DHCP)">Föregående</a><a class="nextlinks-next" href="DPDK.html" title="Data Plane Development Kit">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Time Synchronisation</h1></div>
<div class="region">
<div class="contents">
<p class="para">NTP är ett TCP/IP protokoll för synkronisering av tid över ett nätverk. I grund och botten är det en klient som frågar en server efter nuvarande tid och använder det för att ställa in sin egen klocka.</p>
<p class="para">
Behind this simple description, there is a lot of complexity - there are tiers of NTP servers, with the tier one NTP servers connected to atomic clocks, and tier two and three servers spreading the load of actually handling requests across the Internet. Also the client software is a lot more complex than you might think - it has to factor out communication delays, and adjust the time in a way that does not upset all the other processes that run on the server. But luckily all that complexity is hidden from you! 
</p>
<p class="para">
Ubuntu by default uses <span class="em emphasis">timedatectl / timesyncd</span> to synchronize time and users can optionally use ntpd to serve network time info.
</p>
</div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="NTP.html#timedate-info" title="Synchronizing your systems time">Synchronizing your systems time</a></li>
<li class="links"><a class="xref" href="NTP.html#timeservers" title="Serving NTP">Serving NTP</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-references" title="Referenser">Referenser</a></li>
</ul></div>
<div class="sect2 sect" id="timedate-info"><div class="inner">
<div class="hgroup"><h2 class="title">Synchronizing your systems time</h2></div>
<div class="region">
<div class="contents">
<p class="para">
		Starting with Ubuntu 16.04 <span class="em emphasis">timedatectl / timesyncd</span> (which are part of systemd) replace most of <span class="em emphasis">ntpdate / ntp</span>.
	</p>
<p class="para">
        <span class="app application">timesyncd</span> is available by default and replaces not only <span class="app application">ntpdate</span>, but also the client portion of <span class="app application">ntpd</span>.
		So on top of the one-shot action that <span class="app application">ntpdate</span> provided on boot and network activation, now <span class="app application">timesyncd</span> by default regularly checks and keeps your local time in sync.
		It also stores time updates locally, so that after reboots monotonically advances if applicable.
	</p>
<p class="para">
		If <span class="app application">ntpdate / ntp</span> are installed <span class="app application">timedatectl</span> steps back to let you keep your old setup.
		That shall ensure that no two time syncing services are fighting and also to retain any kind of old behaviour/config that you had through an upgrade.
		But it also implies that on an upgrade from a former release ntp/ntpdate might still be installed and therefore renders the new systemd based services disabled.
	</p>
<p class="para">
		<span class="app application">ntpdate</span> is considered deprecated in favour of <span class="app application">timedatectl</span> and thereby no more installed by default.
	</p>
</div>
<div class="sect3 sect" id="timedate-config"><div class="inner">
<div class="hgroup"><h3 class="title">Configuring timedatectl and timesyncd</h3></div>
<div class="region"><div class="contents">
<p class="para">
		The current status of time and time configuration via <span class="app application">timedatectl</span> and <span class="app application">timesyncd</span> can be checked with <span class="cmd command">timedatectl status</span>.
	</p>
<div class="screen"><pre class="contents ">$ timedatectl status
      Local time: Mo 2017-06-26 12:16:16 CEST
  Universal time: Mo 2017-06-26 10:16:16 UTC
        RTC time: Mo 2017-06-26 10:16:16
       Time zone: Europe/Berlin (CEST, +0200)
 Network time on: yes
NTP synchronized: yes
 RTC in local TZ: no
</pre></div>
<p class="para">
Via <span class="app application">timedatectl</span> an admin can control the timezone, how the system clock should relate to the hwclock and if permanent synronization should be enabled or not.
See <span class="cmd command">man timedatectl</span> for more details.
</p>
<p class="para">
        timesyncd itself is still a normal service, so you can check its status also more in detail via.
<div class="screen"><pre class="contents ">$ systemctl status systemd-timesyncd
. systemd-timesyncd.service - Network Time Synchronization
   Loaded: loaded (/lib/systemd/system/systemd-timesyncd.service; enabled; vendor preset: enabled)
  Drop-In: /lib/systemd/system/systemd-timesyncd.service.d
           |_disable-with-time-daemon.conf
   Active: active (running) since Mo 2017-06-26 11:12:19 CEST; 30min ago
     Docs: man:systemd-timesyncd.service(8)
 Main PID: 12379 (systemd-timesyn)
   Status: "Synchronized to time server [2001:67c:1560:8003::c8]:123 (ntp.ubuntu.com)."
    Tasks: 2
   Memory: 424.0K
      CPU: 12ms
   CGroup: /system.slice/systemd-timesyncd.service
           |_12379 /lib/systemd/systemd-timesyncd

Jun 26 11:12:19 lap systemd[1]: Starting Network Time Synchronization...
Jun 26 11:12:19 lap systemd[1]: Started Network Time Synchronization.
Jun 26 11:12:19 lap systemd-timesyncd[12379]: Synchronized to time server [2001:67c:1560:8003::c8]:123 (ntp.ubuntu.com).
</pre></div>
</p>
<p class="para">
        The nameserver to fetch time for <span class="app application">timedatectl</span> and <span class="app application">timesyncd</span> from can be specified in <span class="file filename">/etc/systemd/timesyncd.conf</span> and additional config files can be stored in <span class="file filename">/etc/systemd/timesyncd.conf.d/</span>.
        The entries for NTP= and FallbackNTP= are space separated lists.
</p>
</div></div>
</div></div>
</div>
</div></div>
<div class="sect2 sect" id="timeservers"><div class="inner">
<div class="hgroup"><h2 class="title">Serving NTP</h2></div>
<div class="region">
<div class="contents"><p class="para">
       If on top of synchronizing your system you also want to serve NTP information you need an ntp server. The most classic and supported one is <span class="app application">ntpd</span>, but it is also very old so there also are <span class="app application">openntpd</span> and <span class="app application">chrony</span> as alternatives available in the archive.
   </p></div>
<div class="sect3 sect" id="ntpd"><div class="inner">
<div class="hgroup"><h3 class="title">ntpd</h3></div>
<div class="region"><div class="contents"><p class="para">
   The ntp daemon ntpd calculates the drift of your system clock and continuously adjusts it, so there are no large corrections that could
   lead to inconsistent logs for instance. The cost is a little processing power and memory, but for a modern server this is negligible.
   </p></div></div>
</div></div>
<div class="sect3 sect" id="ntp-installation"><div class="inner">
<div class="hgroup"><h3 class="title">Installation</h3></div>
<div class="region"><div class="contents">
<p class="para">
   To install ntpd, from a terminal prompt enter:
   </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install ntp</span>
</pre></div>
</div></div>
</div></div>
<div class="sect3 sect" id="timeservers-conf"><div class="inner">
<div class="hgroup"><h3 class="title">Konfiguration</h3></div>
<div class="region"><div class="contents">
<p class="para">
  Edit <span class="file filename">/etc/ntp.conf</span> to add/remove server lines.
  By default these servers are configured:
  </p>
<div class="code"><pre class="contents "># Use servers from the NTP Pool Project. Approved by Ubuntu Technical Board
# on 2011-02-08 (LP: #104525). See http://www.pool.ntp.org/join.html for
# more information.
server 0.ubuntu.pool.ntp.org
server 1.ubuntu.pool.ntp.org
server 2.ubuntu.pool.ntp.org
server 3.ubuntu.pool.ntp.org
</pre></div>
<p class="para">
	  After changing the config file you have to reload the
          <span class="app application">ntpd</span>:
	  </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo systemctl reload ntp.service</span>
</pre></div>
<p class="para">
	   Of the pool number 2.ubuntu.pool.ntp.org as well as ntp.ubuntu.com also support ipv6 if needed.
	   If one needs to force ipv6 there also is ipv6.ntp.ubuntu.com which is not configured by default.
</p>
</div></div>
</div></div>
<div class="sect3 sect" id="ntp-status"><div class="inner">
<div class="hgroup"><h3 class="title">View status</h3></div>
<div class="region"><div class="contents">
<p class="para">
  Use ntpq to see more info: 
  </p>
<div class="screen"><pre class="contents "><span class="cmd command"># sudo ntpq -p</span>
<span class="output computeroutput">     remote           refid      st t when poll reach   delay   offset  jitter
==============================================================================
+stratum2-2.NTP. 129.70.130.70    2 u    5   64  377   68.461  -44.274 110.334
+ntp2.m-online.n 212.18.1.106     2 u    5   64  377   54.629  -27.318  78.882
*145.253.66.170  .DCFa.           1 u   10   64  377   83.607  -30.159  68.343
+stratum2-3.NTP. 129.70.130.70    2 u    5   64  357   68.795  -68.168 104.612
+europium.canoni 193.79.237.14    2 u   63   64  337   81.534  -67.968  92.792</span>
</pre></div>
</div></div>
</div></div>
<div class="sect3 sect" id="ntp-pps"><div class="inner">
<div class="hgroup"><h3 class="title">PPS Support</h3></div>
<div class="region"><div class="contents"><p class="para">
Since 16.04 ntp supports PPS discipline which can be used to augment ntp with local timesources for better accuracy.
For more details on configuration see the external pps ressource listed below.
  </p></div></div>
</div></div>
</div>
</div></div>
<div class="sect2 sect" id="ntp-references"><div class="inner">
<div class="hgroup"><h2 class="title">Referenser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
  	    <p class="para">
          See the <a href="https://help.ubuntu.com/community/UbuntuTime" class="ulink" title="https://help.ubuntu.com/community/UbuntuTime">Ubuntu Time</a> wiki page for more information.
        </p>
      </li>
<li class="list itemizedlist">
  	    <p class="para">
          <a href="http://www.ntp.org/" class="ulink" title="http://www.ntp.org/">ntp.org, home of the Network Time Protocol project</a>
        </p>
      </li>
<li class="list itemizedlist">
  	    <p class="para">
            <a href="https://www.freedesktop.org/software/systemd/man/timedatectl.html" class="ulink" title="https://www.freedesktop.org/software/systemd/man/timedatectl.html">Freedesktop.org info on timedatectl</a>
        </p>
      </li>
<li class="list itemizedlist">
  	    <p class="para">
            <a href="https://www.freedesktop.org/software/systemd/man/systemd-timesyncd.service.html#" class="ulink" title="https://www.freedesktop.org/software/systemd/man/systemd-timesyncd.service.html#">Freedesktop.org info on systemd-timesyncd service</a>
        </p>
      </li>
<li class="list itemizedlist">
  	    <p class="para">
		    <a href="http://www.ntp.org/ntpfaq/NTP-s-config-adv.htm#S-CONFIG-ADV-PPS" class="ulink" title="http://www.ntp.org/ntpfaq/NTP-s-config-adv.htm#S-CONFIG-ADV-PPS">ntp.org faq on configuring PPS</a>
        </p>
      </li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="dhcp.html" title="Dynamic Host Configuration Protocol (DHCP)">Föregående</a><a class="nextlinks-next" href="DPDK.html" title="Data Plane Development Kit">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
