<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Visning och skärm</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 24.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Visning och skärm</span></h1></div>
<div class="region">
<div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="look-resolution.html.sv" title="Ändra skärmens upplösning eller orientering"><span class="title">Ändra skärmens upplösning eller orientering</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra upplösningen på skärmen och dess orientering (rotation).</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="display-dual-monitors.html.sv" title="Anslut en andra skärm till din dator"><span class="title">Anslut en andra skärm till din dator</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in en extra skärm.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="display-night-light.html.sv" title="Justera färgtemperaturen för din skärm"><span class="title">Justera färgtemperaturen för din skärm</span><span class="linkdiv-dash"> — </span><span class="desc">Nattbelysning ändrar färgen på dina skärmar enligt tiden på dygnet.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="display-brightness.html.sv" title="Ställ in ljusstyrka"><span class="title">Ställ in ljusstyrka</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra skärmens ljusstyrka för att göra den läsligare i starkt ljus.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="display-blank.html.sv" title="Ställ in tiden för skärmtömning"><span class="title">Ställ in tiden för skärmtömning</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra tiden till skärmtömning för att spara ström.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="look-background.html.sv" title="Ändra utseendet för ditt skrivbord"><span class="title">Ändra utseendet för ditt skrivbord</span><span class="linkdiv-dash"> — </span><span class="desc">Välj en stil och ställ in en bakgrund.</span></a></div>
</div>
</div></div></div></div></div>
<section id="problems"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Problem</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="session-screenlocks.html.sv" title="Skärmen låser sig själv allt för snabbt"><span class="title">Skärmen låser sig själv allt för snabbt</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra hur länge det tar innan skärmen låser sig själv i <span class="gui">Skärmlås</span>-inställningarna.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="look-display-fuzzy.html.sv" title="Varför ser saker otydliga/pixellerade ut på min skärm?"><span class="title">Varför ser saker otydliga/pixellerade ut på min skärm?</span><span class="linkdiv-dash"> — </span><span class="desc">Skärmupplösningen kan vara felaktigt inställd.</span></a></div>
</div>
<div class="links-divs"><div class="linkdiv "><a class="linkdiv" href="power-whydim.html.sv" title="Varför tonas min skärm ner efter ett tag?"><span class="title">Varför tonas min skärm ner efter ett tag?</span><span class="linkdiv-dash"> — </span><span class="desc">Skärmen tonas ner när datorn är oanvänd för att spara ström.</span></a></div></div>
</div></div></div></div></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — Få GNOME att arbeta för dig, från hårdvarukontroll till sekretessinställningar.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
