<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Trådbunden anslutning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Trådbunden anslutning</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="net-manual.html" title="Ange nätverksinställningar manuellt"><span class="title">Ange nätverksinställningar manuellt</span><span class="linkdiv-dash"> — </span><span class="desc">Om nätverksinställningar inte tilldelas automatiskt kan du behöva mata in dem själv.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-vpn-connect.html" title="Anslut till ett VPN"><span class="title">Anslut till ett VPN</span><span class="linkdiv-dash"> — </span><span class="desc">VPN låter dig ansluta till ett lokalt nätverk via internet. Läs mer om hur du ställer in en VPN-anslutning.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wired-connect.html" title="Anslut till ett trådbundet (Ethernet) nätverk"><span class="title">Anslut till ett trådbundet (Ethernet) nätverk</span><span class="linkdiv-dash"> — </span><span class="desc">För att ställa in de flesta trådbundna anslutningar, är allt du behöver göra att ansluta nätverkskabeln.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-fixed-ip-address.html" title="Skapa en anslutning med en fast IP-adress"><span class="title">Skapa en anslutning med en fast IP-adress</span><span class="linkdiv-dash"> — </span><span class="desc">Med en statisk IP-adress kan det bli enklare att utföra vissa nätverkstjänster från din dator.</span></a></div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a><span class="desc"> — <span class="link"><a href="net-wireless.html" title="Trådlös anslutning">Trådlöst</a></span>, <span class="link"><a href="net-wired.html" title="Trådbunden anslutning">trådbundet</a></span>, <span class="link"><a href="net-problem.html" title="Nätverksproblem">anslutnings-problem</a></span>, <span class="link"><a href="net-browser.html" title="Webbläsare">webbnavigering</a></span>, <span class="link"><a href="net-email.html" title="E-post &amp; e-postmjukvara">e-postkonton</a></span>, <span class="link"><a href="net-chat.html" title="Chatt &amp; sociala medier">snabbmeddelanden</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
