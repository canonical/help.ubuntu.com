<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="600" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-search2.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2">
      <ns0:stop id="stop3964-5-0-1-9-6-6" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68893" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:linearGradient id="linearGradient6868-5-7-5-4-3" ns1:collect="always">
      <ns0:stop id="stop6870-84-7-0-1-8" offset="0" style="stop-color: rgb(0, 0, 0); stop-opacity: 1;"/>
      <ns0:stop id="stop6872-0-5-0-7-1" offset="1" style="stop-color: rgb(0, 0, 0); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68891" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68897" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68895" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68901" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68899" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68905" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68903" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68909" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68907" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68913" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68911" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68917" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68915" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68921" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68919" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68925" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68923" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2-0">
      <ns0:stop id="stop3964-5-0-1-9-6-6-34" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6-4" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7-0"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3-6" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient r="46.177555" fy="152.54469" fx="154.30887" cy="152.54469" cx="154.30887" gradientTransform="matrix(3.8062827,-4.3447397e-8,2.2199035e-8,1.944784,116.22821,273.72246)" gradientUnits="userSpaceOnUse" id="radialGradient25776" ns4:href="#linearGradient5467" ns1:collect="always"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient5467">
      <ns0:stop style="stop-color:#ffffff;stop-opacity:1;" offset="0" id="stop5469"/>
      <ns0:stop style="stop-color:#ffffff;stop-opacity:0.7173913" offset="1" id="stop5471"/>
    </ns0:linearGradient>
    <ns0:radialGradient r="46.177555" fy="152.54469" fx="154.30887" cy="152.54469" cx="154.30887" gradientTransform="matrix(3.8062827,-4.3447397e-8,2.2199035e-8,1.944784,116.22821,273.72246)" gradientUnits="userSpaceOnUse" id="radialGradient25826" ns4:href="#linearGradient5467" ns1:collect="always"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-7">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9-2" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9-2" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6-2" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath987-2-4-1">
      <ns0:circle r="60" cy="236" cx="63.999996" id="circle989-0-6-1" style="display:inline;opacity:1;fill:#3584e4;fill-opacity:1;stroke:none;stroke-width:4.28571415;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="364.52772" ns1:cy="139.55062" ns1:document-units="px" ns1:current-layer="layer2" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="1581" ns1:window-height="1373" ns1:window-x="977" ns1:window-y="27" ns1:window-maximized="0" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0" showguides="true" ns1:guide-bbox="true">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
    <ns2:guide orientation="1,0" position="232,36" id="guide8431" ns1:locked="false"/>
    <ns2:guide orientation="1,0" position="443,51" id="guide8433" ns1:locked="false"/>
    <ns2:guide orientation="1,0" position="178,52" id="guide8535" ns1:locked="false"/>
    <ns2:guide orientation="1,0" position="280,356" id="guide10569" ns1:locked="false"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-892.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="656" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-440)">
    <ns0:g id="g11020" transform="translate(-35,-228.36217)">
      <ns0:path transform="translate(2,453.36217)" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" ns2:ry="17" ns2:rx="17" ns2:cy="278" ns2:cx="120" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
      <ns0:text id="text11016" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan11018" ns2:role="line" style="font-size:14px;line-height:1.25">2</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2.25294995;marker:none;enable-background:new" d="M 118.96098,501.18656 H 720.4075 v 38.66458 c 0,0 -3.02489,-7.96537 -8.33509,-8.23089 l -585.64715,0.79654 c -3.45166,-0.26551 -7.46428,4.13041 -7.46428,4.13041 z" id="rect10989-4" ns1:connector-curvature="0" ns2:nodetypes="ccccccc"/>
    <ns0:rect style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:2.25294995;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:new" id="rect10923-0" width="600.78668" height="450.59" x="119.66641" y="501.62646"/>
    <ns0:path id="path10955-1" style="fill:none;stroke:#000000;stroke-width:1.78223312px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" d="m 719.85155,539.75089 c 0,-4.42934 -3.59068,-8.02005 -8.02006,-8.02005 H 127.56697 c -4.42936,0 -8.02005,3.59071 -8.02005,8.02005" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:9.01179981px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.75098336" x="419.94446" y="522.79474" id="text10972-5"><ns0:tspan ns2:role="line" id="tspan10974-5" x="419.94446" y="522.79474" style="font-size:15.96732807px;line-height:1.25;stroke-width:0.75098336">14:30</ns0:tspan></ns0:text>
    <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 225.94527,530.22888 h -97.62731 c -4.42937,0 -8.02005,3.5907 -8.02005,8.02005" style="fill:none;stroke:#000000;stroke-width:3.75491667;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" id="path17186"/>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:9.01179981px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.75098336" x="126.4698" y="522.79474" id="text56758"><ns0:tspan ns2:role="line" id="tspan56760" x="126.4698" y="522.79474" style="font-size:15.96732807px;line-height:1.25;stroke-width:0.75098336">Aktiviteter</ns0:tspan></ns0:text>
    <ns0:g style="display:inline" ns1:label="audio-volume-medium" transform="translate(640.40993,291.45883)" id="g5525">
      <ns0:path ns1:connector-curvature="0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none" d="m 20,222 h 2.484375 L 25.453129,219 26,219.0156 v 11 l -0.475297,8.3e-4 L 22.484375,227 H 20 Z" id="path5533" ns2:nodetypes="ccccccccc"/>
      <ns0:rect ns1:label="audio-volume-high" y="217" x="20" height="16" width="16" id="rect5535" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none"/>
      <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3718-5" style="display:inline;fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:type="arc" clip-path="url(#clipPath6279-7-9-7)"/>
      <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" ns2:type="arc" style="display:inline;fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" id="path3726-1" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" clip-path="url(#clipPath6265-3-4-4)"/>
      <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3728-0" style="display:inline;opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:type="arc" clip-path="url(#clipPath6259-8-81-2)"/>
    </ns0:g>
    <ns0:g style="display:inline" id="g4692-3" ns1:label="system-shutdown" transform="translate(640.40993,-179.54117)">
      <ns0:rect width="16" height="16" rx="0.14408804" ry="0.15129246" x="40" y="688" id="rect10837-3-0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none;enable-background:new"/>
      <ns0:path ns2:type="arc" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" id="path3869-2" ns2:cx="48" ns2:cy="696" ns2:rx="7" ns2:ry="7" d="m 51.52343,689.95141 a 7,7 0 0 1 3.233191,7.87837 7,7 0 0 1 -6.766907,5.17021 7,7 0 0 1 -6.751683,-5.19008 7,7 0 0 1 3.25633,-7.86883" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" ns2:start="5.239857" ns2:end="4.1878597" ns2:open="true"/>
      <ns0:path ns1:connector-curvature="0" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="m 48,689 v 5" id="path4710" ns2:nodetypes="cc"/>
    </ns0:g>
    <ns0:g style="display:inline" ns1:label="network-wired" transform="translate(617.48279,292.54116)" id="g12661">
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" id="rect12673" width="16" height="16" x="20" y="217" ns1:label="audio-volume-high"/>
      <ns0:path ns1:connector-curvature="0" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:Sans;-inkscape-font-specification:Sans;text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;baseline-shift:baseline;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;enable-background:accumulate" d="m -55.25,-40 c -0.952203,0 -1.75,0.7978 -1.75,1.75 v 4.5 c 0,0.9522 0.797797,1.75 1.75,1.75 h 0.125 l -0.78125,1.5625 L -56.625,-29 h 1.625 6 1.625 L -48.09375,-30.4375 -48.875,-32 h 0.125 c 0.952203,0 1.75,-0.7978 1.75,-1.75 v -4.5 c 0,-0.9522 -0.797797,-1.75 -1.75,-1.75 z m 0.25,2 h 6 v 4 h -6 z" transform="translate(80,257)" id="rect12675"/>
      <ns0:path ns1:connector-curvature="0" transform="translate(-60.0003,30)" id="path12679" d="m 88,196 v 4" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
      <ns0:path ns1:connector-curvature="0" id="path12681" d="m 21.99975,231 h 12" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
    </ns0:g>
    <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:3;marker:none;enable-background:accumulate" d="m 710.51717,516.87513 -3.74999,3.75 -3.75001,-3.75 z" id="rect12003" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
    <ns0:g id="g11578" transform="matrix(1.256737,0,0,1.256737,695.80575,-123.70167)">
      <ns0:g style="display:inline;stroke-width:0.93333334;enable-background:new" transform="matrix(0.09738145,0,0,0.09738145,-215.1,597.27741)" id="g912-6">
        <ns0:circle r="224" cy="43.999989" cx="256" id="circle1036" style="display:inline;opacity:1;fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:14.9333334;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="ccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccc" ns1:connector-curvature="0" id="path991" d="m 38,176 v 4 l 10,8 v 8 l 8,8 h 4 v -4 l 6,-6 v -4 l 4,-4 v -10 z m -4,16 H 4 c 0,0 0.5090211,40.4419 0,40 l 20,18 v -6 l -4,-4 6,-6 h 4 l 4,4 0.12494,-8.4018 L 40,224 h 4 v -4 l 4,-4 v -6 L 43.727619,206.12499 34,206 v 8 h -4 l -4,-4 v -4 l 6,-6 h 6 v -4 z m 60,2 -6,6 v 4 h 6 v -2.14287 h 4 v 4.26786 L 96,208 H 86 v 4 h -4 v 6 h -8 v 8 h 10 v -4 h 8 v 2 l 4,4 h 2 v -2 l -2,-2 v -2 h 4 l 6,6 h 6 v 2 l -2,2 h -4 l 18,18 V 194 H 96 Z m 12,38 H 94 l -2,-2 H 78 l -8,8 v 8 l 8,8 h 6 l 4,4 v 2 l 2,2 v 12 l 14,14 h 8 v -30 l 4,-4 v -8 l -10,-10 z m -2,-12 h 4 l 6,6 h -4 z m -74,28 -4,4 v 10 l 8.12494,8.14285 L 34,296 h 8 v -8 l 6,-6 v -4 l 6,-6 v -4 l 4,-4 v -8 l -4,-4 h -8 l -4,-4 z" clip-path="url(#clipPath987-2-4-1)" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.01129821px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:accumulate" transform="matrix(0.3507037,0,0,0.3507037,-212.61539,518.79611)"/>
      <ns0:g transform="matrix(0.12007553,0,0,0.12007553,-302.36423,551.40018)" id="g6008" style="display:inline;opacity:1;stroke:#000000;enable-background:new">
        <ns0:circle r="36.270779" cy="372.21783" cx="883.60425" id="path3066-4" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:16.92636299;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
        <ns0:circle r="68.971695" cy="372.2179" cx="883.60431" id="path3941-2" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:11.69271851;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
        <ns0:circle r="103.1213" cy="372.21796" cx="883.60437" id="path3943-0" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:5.99500418;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
      </ns0:g>
      <ns0:g transform="matrix(0.3635574,0,0,0.3635574,-213.43802,520.12533)" id="g6092" style="display:inline;enable-background:new">
        <ns0:g id="g6087">
          <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:new" ns2:nodetypes="cccssccc" id="path3970-7-4" d="m 47.589745,209.314 -47.7665216,46.36163 21.7759096,0.70244 c 0,0 -9.131831,18.96611 -9.131831,18.96611 -2.8097966,8.42939 9.834282,11.59041 11.941628,5.26838 0,0 8.42939,-18.96612 8.42939,-18.96612 l 15.453872,16.50755 z" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g11589">
      <ns0:path ns1:connector-curvature="0" id="path1558" d="m -206.74531,640.32202 a 4.3626888,4.3626888 0 0 0 -4.36271,4.36268 4.3626888,4.3626888 0 0 0 2.90847,4.10778 v 23.77753 a 4.3626888,4.3626888 0 0 0 -2.90847,4.10777 4.3626888,4.3626888 0 0 0 4.36271,4.36272 4.3626888,4.3626888 0 0 0 3.77403,-2.18138 h 24.4471 a 4.3626888,4.3626888 0 0 0 3.77188,2.18138 4.3626888,4.3626888 0 0 0 4.36273,-4.36272 4.3626888,4.3626888 0 0 0 -2.90849,-4.10777 v -23.77753 a 4.3626888,4.3626888 0 0 0 2.90849,-4.10778 4.3626888,4.3626888 0 0 0 -4.36273,-4.36268 4.3626888,4.3626888 0 0 0 -4.29664,3.63558 h -23.39546 a 4.3626888,4.3626888 0 0 0 -4.30091,-3.63558 z m 3.77403,6.54404 h 24.4471 a 4.3626888,4.3626888 0 0 0 0.0953,0.16622 l -3.76978,3.76979 a 2.9084593,2.9084593 0 0 0 -1.27883,-0.30046 2.9084593,2.9084593 0 0 0 -2.81192,2.18131 h -8.91635 a 2.9084593,2.9084593 0 0 0 -2.81403,-2.18131 2.9084593,2.9084593 0 0 0 -1.28025,0.2989 l -3.77121,-3.77122 a 4.3626888,4.3626888 0 0 0 0.10021,-0.1635 z m -2.31981,2.05637 4.36835,4.36838 a 2.9084593,2.9084593 0 0 0 -0.004,0.11939 2.9084593,2.9084593 0 0 0 1.45422,2.51577 v 9.51216 a 2.9084593,2.9084593 0 0 0 -1.45422,2.51438 2.9084593,2.9084593 0 0 0 0.2989,1.28026 l -3.77118,3.7712 a 4.3626888,4.3626888 0 0 0 -0.89044,-0.43385 z m 29.08458,0 v 23.64758 a 4.3626888,4.3626888 0 0 0 -0.89326,0.431 l -3.76977,-3.7698 a 2.9084593,2.9084593 0 0 0 0.30046,-1.2788 2.9084593,2.9084593 0 0 0 -1.45421,-2.51583 v -9.51211 a 2.9084593,2.9084593 0 0 0 1.45421,-2.51437 2.9084593,2.9084593 0 0 0 -0.004,-0.12056 z m -19.89481,6.66903 h 10.70365 a 2.9084593,2.9084593 0 0 0 0.46579,0.33441 v 9.51216 a 2.9084593,2.9084593 0 0 0 -1.35768,1.78723 h -8.91638 a 2.9084593,2.9084593 0 0 0 -1.35979,-1.78868 v -9.51211 a 2.9084593,2.9084593 0 0 0 0.46441,-0.33285 z m 0,14.54226 h 10.70365 a 2.9084593,2.9084593 0 0 0 1.92003,0.72713 2.9084593,2.9084593 0 0 0 0.12055,-0.004 l 4.46211,4.46211 a 4.3626888,4.3626888 0 0 0 -0.15413,0.63199 h -23.39546 a 4.3626888,4.3626888 0 0 0 -0.16038,-0.62985 l 4.46567,-4.46564 a 2.9084593,2.9084593 0 0 0 0.11939,0.004 2.9084593,2.9084593 0 0 0 1.91862,-0.72715 z" style="color:#000000;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:sans-serif;font-variant-ligatures:normal;font-variant-position:normal;font-variant-caps:normal;font-variant-numeric:normal;font-variant-alternates:normal;font-feature-settings:normal;text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;text-decoration-style:solid;text-decoration-color:#000000;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-orientation:mixed;dominant-baseline:auto;baseline-shift:baseline;text-anchor:start;white-space:normal;shape-padding:0;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2.90845919;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:new"/>
    </ns0:g>
    <ns0:g id="g11597" transform="matrix(0.7698253,0,0,0.7698253,340.83868,259.65604)">
      <ns0:rect ry="3.1104455" rx="3.1104455" y="696.49127" x="-207.98987" height="41.991028" width="34.21489" id="rect15435-6" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:1.45422959;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:path style="display:inline;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.00433091px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" d="m -203.97049,698.99079 c -0.80564,0 -1.45422,0.64858 -1.45422,1.45423 v 10.49772 h 29.08459 v -10.49772 c 0,-0.80565 -0.64859,-1.45423 -1.45423,-1.45423 z m -1.45422,12.67906 v 10.90672 h 29.08459 v -10.90672 z m 0,11.63384 v 10.54316 c 0,0.80565 0.64858,1.45423 1.45422,1.45423 h 26.17614 c 0.80564,0 1.45423,-0.64858 1.45423,-1.45423 v -10.54316 z" id="rect15441-8" ns1:connector-curvature="0" ns2:nodetypes="ssccsssccccccsssscc"/>
      <ns0:g transform="matrix(0.3635574,0,0,0.3635574,-214.15009,632.41434)" id="g1088">
        <ns0:path style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.01184966px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" d="m 552,443 c -1.662,0 -3,1.338 -3,3 v 4 1 h 4 0.0312 l -0.0156,-2 H 569 v 2 H 569.0312 573 v -1 -4 c 0,-2 -1.338,-3 -3,-3 z" transform="translate(-497,-247)" id="path26035" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:use height="100%" width="100%" transform="translate(8.4388398e-7,11.633826)" id="use1090" ns4:href="#g1088" y="0" x="0"/>
      <ns0:use x="0" y="0" ns4:href="#g1088" id="use1092" transform="translate(8.4388398e-7,23.267663)" width="100%" height="100%"/>
    </ns0:g>
    <ns0:g id="g11604">
      <ns0:path ns1:connector-curvature="0" id="rect854" d="m -207.12029,754.15227 c -1.70883,0 -3.08454,1.3757 -3.08454,3.08454 v 3.85565 26.98973 3.08454 c 0,1.70883 1.37571,3.08454 3.08454,3.08454 h 33.92993 c 1.70883,0 3.08453,-1.37571 3.08453,-3.08454 v -3.08454 -26.98973 -3.85565 c 0,-1.70884 -1.3757,-3.08454 -3.08453,-3.08454 z" style="display:inline;opacity:1;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:1.45422959;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
      <ns0:rect style="display:inline;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.00407583px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" id="rect858" width="34.901512" height="31.99304" x="-207.60608" y="-788.74408" rx="1.4542296" ry="1.4542185" transform="scale(1,-1)"/>
      <ns0:g style="display:inline;fill:#ffffff;enable-background:new" transform="matrix(0.3635574,0,0,0.3635574,-214.15012,687.6751)" id="g866">
        <ns0:path ns1:connector-curvature="0" id="path862" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:medium;line-height:1.25;font-family:'Source Code Pro';-inkscape-font-specification:'Source Code Pro, Bold';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.24999999" d="M 44.012301,210.88755 30,203.27182 V 208 l 9.710724,4.62951 v 0.1422 L 30,218 v 4.72818 l 14.012301,-8.21451 z" ns2:nodetypes="ccccccccc"/>
        <ns0:path ns2:nodetypes="ccccc" ns1:connector-curvature="0" id="path864" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:medium;line-height:1.25;font-family:'Source Code Pro';-inkscape-font-specification:'Source Code Pro, Bold';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.24999999" d="m 47.999998,226 2e-6,4 h 16.00001 l -2e-6,-4 z"/>
      </ns0:g>
    </ns0:g>
    <ns0:rect style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:2.25294995;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:new" id="rect11062-3" width="218.1161" height="36.352684" x="306.49579" y="549.53668" rx="18.176342" ry="18.176342"/>
    <ns0:ellipse cy="565.49219" cx="500.47089" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:3.03790092;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" id="path27918" rx="6.8430524" ry="6.8352771"/>
    <ns0:path ns1:connector-curvature="0" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:3.03790092;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" d="m 505.79327,570.8085 6.08271,6.0758" id="path27941" ns2:nodetypes="cc"/>
    <ns0:rect y="555.61896" x="490.58646" height="24.303207" width="24.303211" id="rect1431" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.70638272;fill:none;stroke:none;stroke-width:1.50196671;marker:none;enable-background:accumulate"/>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="323.60797" y="571.51361" id="text57298"><ns0:tspan ns2:role="line" id="tspan57300" x="323.60797" y="571.51361" style="font-size:14px;line-height:1.25">kon</ns0:tspan></ns0:text>
    <ns0:text id="text8415" y="902.51361" x="232.60797" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="902.51361" x="232.60797" id="tspan8417" ns2:role="line" style="font-size:12px;line-height:1.25">Konton</ns0:tspan></ns0:text>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="232.60797" y="922.51361" id="text8419"><ns0:tspan ns2:role="line" id="tspan8421" x="232.60797" y="922.51361" style="font-size:12px;line-height:1.25">https://accounts.google.com/ServiceLogin?service=oz&amp;con...</ns0:tspan></ns0:text>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="281.60797" y="817.51361" id="text8423"><ns0:tspan ns2:role="line" id="tspan8425" x="281.60797" y="817.51361" style="font-size:12px;line-height:1.25">konfiguration</ns0:tspan></ns0:text>
    <ns0:text id="text8427" y="859.51361" x="281.60797" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="859.51361" x="281.60797" id="tspan8429" ns2:role="line" style="font-size:12px;line-height:1.25">fontconfig</ns0:tspan></ns0:text>
    <ns0:text id="text8435" y="817.51361" x="482" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="817.51361" x="482" id="tspan8437" ns2:role="line" style="font-size:12px;line-height:1.25">system-config-http.zip</ns0:tspan></ns0:text>
    <ns0:text id="text8457" y="724.51361" x="280.60797" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="724.51361" x="280.60797" id="tspan8459" ns2:role="line" style="font-size:12px;line-height:1.25">Ikonriktlinjer</ns0:tspan></ns0:text>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="280.60797" y="759.51361" id="text8461"><ns0:tspan ns2:role="line" id="tspan8463" x="280.60797" y="759.51361" style="font-size:12px;line-height:1.25">fontconfig</ns0:tspan></ns0:text>
    <ns0:rect style="color:#000000;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect10535" width="30" height="28" x="232" y="707"/>
    <ns0:rect y="742" x="232" height="28" width="30" id="rect10537" style="color:#000000;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:g id="g7262" ns1:label="package-x-generic" transform="matrix(2,0,0,2,346.9996,-3)">
      <ns0:rect y="398" x="48" height="16" width="16" id="rect7264" style="opacity:0.51464431;color:#bebebe;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 51.0002,406 10,0 0,7.05898 c 0,0.4922 -0.47266,0.9375 -0.99609,0.9375 l -8.00391,0 C 51.46114,413.99648 51.0002,413.56684 51.0002,412.99648 Z" id="rect7268" ns1:connector-curvature="0" ns2:nodetypes="ccccccc"/>
      <ns0:path style="fill:none;stroke:#bebebe;stroke-width:2;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 52.0002,406.4375 0,-1 2.815996,-3.45781" id="path7270" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
      <ns0:path style="fill:none;stroke:#bebebe;stroke-width:2;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 60.03145,406.5 0,-1 -2.99798,-0.5243" id="path7272" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
    </ns0:g>
    <ns0:g id="g4958" ns1:label="folder" transform="matrix(1.9999998,0,0,1.9999998,-183.99956,-1196.9998)" style="display:inline">
      <ns0:path ns2:nodetypes="ccccccccccsccccccccccc" id="rect3845" d="m 208.53105,997 c -0.28913,0 -0.53125,0.24212 -0.53125,0.53125 l 0,13.93755 c 0,0.2985 0.23264,0.5312 0.53125,0.5312 l 14.9375,0 c 0.2986,0 0.53125,-0.2326 0.53125,-0.5312 l 0,-8.9376 c 0,-0.2891 -0.24212,-0.5312 -0.53125,-0.5312 l -12.46875,0 0,7.5 c 0,0.277 -0.223,0.5 -0.5,0.5 -0.277,0 -0.5,-0.223 -0.5,-0.5 l 0,-8 c 0,-0.277 0.223,-0.5 0.5,-0.5 l 2.96875,0 8.53125,0 0,-1.4062 c 0,-0.3272 -0.26666,-0.5938 -0.59375,-0.5938 l -7.40625,0 0,-1.46875 C 213.9998,997.2421 213.75768,997 213.46855,997 Z" style="fill:#bebebe;fill-opacity:1;stroke:none;display:inline" ns1:connector-curvature="0"/>
      <ns0:rect y="996" x="207.9998" height="16" width="16" id="rect14152" style="color:#bebebe;fill:none;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:g>
    <ns0:g style="display:inline" transform="matrix(1.9999998,0,0,1.9999998,-183.99956,-1156.9998)" ns1:label="folder" id="g10595">
      <ns0:path ns1:connector-curvature="0" style="fill:#bebebe;fill-opacity:1;stroke:none;display:inline" d="m 208.53105,997 c -0.28913,0 -0.53125,0.24212 -0.53125,0.53125 l 0,13.93755 c 0,0.2985 0.23264,0.5312 0.53125,0.5312 l 14.9375,0 c 0.2986,0 0.53125,-0.2326 0.53125,-0.5312 l 0,-8.9376 c 0,-0.2891 -0.24212,-0.5312 -0.53125,-0.5312 l -12.46875,0 0,7.5 c 0,0.277 -0.223,0.5 -0.5,0.5 -0.277,0 -0.5,-0.223 -0.5,-0.5 l 0,-8 c 0,-0.277 0.223,-0.5 0.5,-0.5 l 2.96875,0 8.53125,0 0,-1.4062 c 0,-0.3272 -0.26666,-0.5938 -0.59375,-0.5938 l -7.40625,0 0,-1.46875 C 213.9998,997.2421 213.75768,997 213.46855,997 Z" id="path10597" ns2:nodetypes="ccccccccccsccccccccccc"/>
      <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect10599" width="16" height="16" x="207.9998" y="996"/>
    </ns0:g>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="491.60797" y="724.51361" id="text10601"><ns0:tspan ns2:role="line" id="tspan10603" x="491.60797" y="724.51361" style="font-size:12px;line-height:1.25">Säkra Linux-behållare</ns0:tspan></ns0:text>
    <ns0:text id="text10605" y="759.51361" x="491.60797" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="759.51361" x="491.60797" id="tspan10607" ns2:role="line" style="font-size:12px;line-height:1.25">Utvecklarkonferens 2012</ns0:tspan></ns0:text>
    <ns0:rect y="707" x="443" height="28" width="30" id="rect10609" style="color:#000000;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:rect style="color:#000000;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect10611" width="30" height="28" x="443" y="742"/>
    <ns0:g transform="matrix(0.5,0,0,0.5,-107.5,363.31891)" id="g24776" ns1:label="documents">
      <ns0:path style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:7;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero" d="m 608.17584,693.39936 -29.90154,9.20048 9.20047,28.43782 L 617.1672,721.83719 Z" id="path24774" ns1:connector-curvature="0"/>
      <ns0:rect y="687.36218" x="573" height="64" width="64" id="rect24747" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:path ns2:nodetypes="cccccc" ns1:connector-curvature="0" id="path21570" d="m 590.85066,695.9724 0,48.284 39.75057,0 0,-39.53456 L 621.52773,695.9724 Z" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:5;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:path ns1:connector-curvature="0" id="path24751" d="m 609.19489,730.79208 11.94524,-1.63633 -3.09102,-20.75399 m -12.80011,-8.22934 -19.02884,2.84563 4.39113,30.31973" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero" ns2:nodetypes="cccccc"/>
      <ns0:path ns1:connector-curvature="0" id="path24749" d="m 608.17584,693.39936 -29.90154,9.20048 9.20047,28.43782 L 617.1672,721.83719 Z" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:path style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:none;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero" d="m 598.29097,704.40685 0,12.82105 -2.46912,2.89508 -2.82186,-3.30866 0,-26.05569 7.05464,0 0,4.5494" id="path24783" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:g transform="translate(-324.07727,68.659424)" id="g25797">
      <ns0:rect y="530.34058" x="673.07727" height="64" width="64" id="rect25795" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:rect ry="2.4805617" rx="2.4805617" y="539.61224" x="717.70361" height="15.50351" width="10.852457" id="rect25714" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:#edf3fb;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:rect ry="2.4805617" rx="2.4805617" y="552.41345" x="718.67584" height="15.193439" width="11.782667" id="rect25716" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:#edf3fb;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:rect ry="2.277133" rx="2.488415" y="565.36646" x="716.48029" height="16.793856" width="15.863646" id="rect25718" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:#edf3fb;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:rect ry="2.4960177" rx="2.4805617" y="534.2077" x="678.05804" height="57.096397" width="48.060883" id="rect25712" style="color:#000000;color-interpolation:sRGB;color-interpolation-filters:linearRGB;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:4;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;clip-rule:nonzero"/>
      <ns0:path style="font-size:23.55376053px;font-style:normal;font-weight:normal;fill:url(#radialGradient25826);fill-opacity:1;stroke:none;display:inline;enable-background:new;font-family:Bitstream Vera Sans" id="path5099" d="m 700.43477,563.41392 c -2e-5,1.41414 0.28918,2.52934 0.86758,3.34562 0.5895,0.81629 1.38479,1.22443 2.38587,1.22443 0.98992,0 1.77964,-0.40814 2.36918,-1.22443 0.58949,-0.82777 0.88425,-1.94298 0.88427,-3.34562 -2e-5,-1.39112 -0.30034,-2.48908 -0.90096,-3.29388 -0.58953,-0.81627 -1.38482,-1.22442 -2.38586,-1.22443 -0.97883,10e-6 -1.763,0.40816 -2.3525,1.22443 -0.5784,0.8048 -0.8676,1.90276 -0.86758,3.29388 m 6.84059,5.19088 c -0.33371,0.81629 -0.87317,1.45437 -1.61839,1.91425 -0.73413,0.44838 -1.59615,0.67258 -2.58607,0.67258 -1.91316,0 -3.47037,-0.71282 -4.67162,-2.13844 -1.19017,-1.43712 -1.78524,-3.30538 -1.78523,-5.60478 -10e-6,-2.29938 0.60062,-4.16764 1.80191,-5.60477 1.20126,-1.43711 2.7529,-2.15567 4.65494,-2.15569 0.98992,2e-5 1.85194,0.22996 2.58607,0.68982 0.74522,0.4599 1.28468,1.09798 1.61839,1.91425 l 0,-2.25916 3.48703,0 0,11.95111 c 1.37922,-0.21844 2.4637,-0.90251 3.25345,-2.05221 0.7897,-1.16119 1.18456,-2.6443 1.18459,-4.44933 -3e-5,-1.14969 -0.16131,-2.22465 -0.48385,-3.2249 -0.32259,-1.01172 -0.81199,-1.93723 -1.46822,-2.77652 -1.0567,-1.40262 -2.38033,-2.48333 -3.97088,-3.24215 -1.57947,-0.75878 -3.2924,-1.13818 -5.13878,-1.1382 -1.29028,2e-5 -2.52492,0.17823 -3.70393,0.53461 -1.17904,0.34493 -2.26909,0.85655 -3.27014,1.53485 -1.6462,1.12672 -2.93089,2.58683 -3.85408,4.38034 -0.91209,1.78205 -1.36813,3.71354 -1.36812,5.79448 -10e-6,1.71306 0.29475,3.32263 0.88427,4.82873 0.60063,1.49461 1.46265,2.81676 2.58608,3.96645 1.11228,1.12671 2.38585,1.98323 3.82071,2.56958 1.44597,0.59784 2.98649,0.89676 4.62157,0.89676 1.40147,0 2.80296,-0.27018 4.20446,-0.81053 1.40147,-0.54036 2.59718,-1.27042 3.58714,-2.19018 l 1.78523,2.79377 c -1.39039,1.1152 -2.90867,1.96598 -4.55484,2.55233 -1.63508,0.59783 -3.29796,0.89675 -4.98862,0.89676 -2.05775,-10e-6 -3.9987,-0.37941 -5.82284,-1.1382 -1.82417,-0.74731 -3.44811,-1.83952 -4.87184,-3.27664 -1.42373,-1.43712 -2.50822,-3.09843 -3.25345,-4.98394 -0.74523,-1.89699 -1.11785,-3.93196 -1.11785,-6.10489 0,-2.09244 0.37818,-4.08716 1.13454,-5.98418 0.75635,-1.89698 1.83527,-3.56404 3.23676,-5.00118 1.40148,-1.42561 3.03098,-2.52931 4.88852,-3.31113 1.86864,-0.78177 3.80402,-1.17266 5.80616,-1.17269 2.49151,3e-5 4.75502,0.49439 6.79053,1.48311 2.03547,0.97726 3.73728,2.39139 5.10542,4.24238 0.83419,1.12673 1.46264,2.35115 1.88534,3.67328 0.43376,1.31067 0.65066,2.69031 0.65069,4.13892 -3e-5,3.11569 -0.90655,5.5358 -2.71955,7.26034 -1.81307,1.72454 -4.37133,2.58682 -7.67481,2.58682 l -0.65069,0 0,-2.65581" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none" x="376.60797" y="675.51361" id="text25881"><ns0:tspan ns2:role="line" id="tspan25883" x="376.60797" y="675.51361" style="font-size:12.00000095px;line-height:1.25">Kontakter</ns0:tspan></ns0:text>
    <ns0:text id="text25885" y="675.51361" x="455.60797" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="675.51361" x="455.60797" id="tspan25887" ns2:role="line" style="font-size:12.00000095px;line-height:1.25">Webb</ns0:tspan></ns0:text>
    <ns0:g transform="matrix(0.65768384,0,0,0.65768384,319.65778,512.94284)" id="g11626">
      <ns0:g id="g11608" transform="matrix(0.09738145,0,0,0.09738145,-215.1,597.27741)" style="display:inline;stroke-width:0.93333334;enable-background:new">
        <ns0:circle style="display:inline;opacity:1;fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:14.9333334;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" id="circle11606" cx="256" cy="43.999989" r="224"/>
      </ns0:g>
      <ns0:path transform="matrix(0.3507037,0,0,0.3507037,-212.61539,518.79611)" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.01129821px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:accumulate" clip-path="url(#clipPath987-2-4-1)" d="m 38,176 v 4 l 10,8 v 8 l 8,8 h 4 v -4 l 6,-6 v -4 l 4,-4 v -10 z m -4,16 H 4 c 0,0 0.5090211,40.4419 0,40 l 20,18 v -6 l -4,-4 6,-6 h 4 l 4,4 0.12494,-8.4018 L 40,224 h 4 v -4 l 4,-4 v -6 L 43.727619,206.12499 34,206 v 8 h -4 l -4,-4 v -4 l 6,-6 h 6 v -4 z m 60,2 -6,6 v 4 h 6 v -2.14287 h 4 v 4.26786 L 96,208 H 86 v 4 h -4 v 6 h -8 v 8 h 10 v -4 h 8 v 2 l 4,4 h 2 v -2 l -2,-2 v -2 h 4 l 6,6 h 6 v 2 l -2,2 h -4 l 18,18 V 194 H 96 Z m 12,38 H 94 l -2,-2 H 78 l -8,8 v 8 l 8,8 h 6 l 4,4 v 2 l 2,2 v 12 l 14,14 h 8 v -30 l 4,-4 v -8 l -10,-10 z m -2,-12 h 4 l 6,6 h -4 z m -74,28 -4,4 v 10 l 8.12494,8.14285 L 34,296 h 8 v -8 l 6,-6 v -4 l 6,-6 v -4 l 4,-4 v -8 l -4,-4 h -8 l -4,-4 z" id="path11610" ns1:connector-curvature="0" ns2:nodetypes="ccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccc"/>
      <ns0:g style="display:inline;opacity:1;stroke:#000000;enable-background:new" id="g11618" transform="matrix(0.12007553,0,0,0.12007553,-302.36423,551.40018)">
        <ns0:circle style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:16.92636299;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none" id="circle11612" cx="883.60425" cy="372.21783" r="36.270779"/>
        <ns0:circle style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:11.69271851;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none" id="circle11614" cx="883.60431" cy="372.2179" r="68.971695"/>
        <ns0:circle style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:5.99500418;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none" id="circle11616" cx="883.60437" cy="372.21796" r="103.1213"/>
      </ns0:g>
      <ns0:g style="display:inline;enable-background:new" id="g11624" transform="matrix(0.3635574,0,0,0.3635574,-213.43802,520.12533)">
        <ns0:g id="g11622">
          <ns0:path ns1:connector-curvature="0" d="m 47.589745,209.314 -47.7665216,46.36163 21.7759096,0.70244 c 0,0 -9.131831,18.96611 -9.131831,18.96611 -2.8097966,8.42939 9.834282,11.59041 11.941628,5.26838 0,0 8.42939,-18.96612 8.42939,-18.96612 l 15.453872,16.50755 z" id="path11620" ns2:nodetypes="cccssccc" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:new"/>
        </ns0:g>
      </ns0:g>
    </ns0:g>
  </ns0:g>
</ns0:svg>
