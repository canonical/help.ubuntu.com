<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>OpenSSH-server</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="remote-administration.html" title="Fjärradministration">Fjärradministration</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="remote-administration.html" title="Fjärradministration">Föregående</a><a class="nextlinks-next" href="puppet.html" title="Puppet">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">OpenSSH-server</h1></div>
<div class="region">
<div class="contents"></div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="openssh-server.html#openssh-introduction" title="Inledning">Inledning</a></li>
<li class="links"><a class="xref" href="openssh-server.html#openssh-installation" title="Installation">Installation</a></li>
<li class="links"><a class="xref" href="openssh-server.html#openssh-configuration" title="Konfiguration">Konfiguration</a></li>
<li class="links"><a class="xref" href="openssh-server.html#openssh-keys" title="SSH-nycklar">SSH-nycklar</a></li>
<li class="links"><a class="xref" href="openssh-server.html#openssh-references" title="Referenser">Referenser</a></li>
</ul></div>
<div class="sect2 sect" id="openssh-introduction"><div class="inner">
<div class="hgroup"><h2 class="title">Inledning</h2></div>
<div class="region"><div class="contents">
<p class="para">
            This section of the Ubuntu Server Guide introduces a powerful collection of tools
            for the remote control of, and transfer of data between, networked computers called <span class="em emphasis">OpenSSH</span>. You will also learn
            about some of the configuration settings possible with the OpenSSH server application and how to change them on your Ubuntu system.
          </p>
<p class="para">
            OpenSSH is a freely available version of the Secure Shell (SSH) protocol family of
            tools for remotely controlling, or transferring files between, computers.
            Traditional tools used to accomplish these functions, such as
	    <span class="app application">telnet</span> or <span class="app application">rcp</span>, are insecure
	    and transmit the user's password in cleartext when used. OpenSSH provides a server
	    daemon and client tools to facilitate secure, encrypted remote control and file
	    transfer operations, effectively replacing the legacy tools.
          </p>
<p class="para">Serverkomponenten i OpenSSH, <span class="app application">sshd</span>, lyssnar kontinuerligt efter klientanslutningar från något av klientverktygen. När en anslutningsförfrågan anländer skapar <span class="app application">sshd</span> korrekt anslutning beroende på vilket klientverktyg som ansluter. Till exempel, om fjärrdatorn ansluter med klientprogrammet <span class="app application">ssh</span> kommer OpenSSH-servern att skapa en fjärrstyrningssession efter att klienten autentiserat sig. Om fjärrdatorn ansluter till OpenSSH-servern med <span class="app application">scp</span> skapar OpenSSH-servern istället en anslutning för säker kopiering av filer mellan servern och klienten efter att klienten autentiserat sig. OpenSSH kan använda flera autentiseringsmetoder, inklusive vanliga lösenord, publik nyckel och <span class="app application">Kerberos</span>-certifikat.</p>
</div></div>
</div></div>
<div class="sect2 sect" id="openssh-installation"><div class="inner">
<div class="hgroup"><h2 class="title">Installation</h2></div>
<div class="region"><div class="contents">
<p class="para">Installationen av OpenSSH-klienten och -servern är enkel. För att installera OpenSSH-klienten på din Ubuntu-dator, kör det här kommandot från en terminalprompt:</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install openssh-client</span>
</pre></div>
<p class="para">För att installera OpenSSH-servern, och relaterade stödfiler, använd det här kommandot från en terminalprompt:</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install openssh-server</span>
</pre></div>
<p class="para">Paketet <span class="app application">openssh-server</span> kan också väljas för installation under installationsprocessen av Server Edition.</p>
</div></div>
</div></div>
<div class="sect2 sect" id="openssh-configuration"><div class="inner">
<div class="hgroup"><h2 class="title">Konfiguration</h2></div>
<div class="region"><div class="contents">
<p class="para">Du kan konfigurera standardbeteendet för OpenSSH-servern <span class="app application">sshd</span>, genom att ändra i filen <span class="file filename">/etc/ssh/sshd_config</span>. För information om konfigurationsmöjligheterna som används i den här filen, kan du med följande kommando, som du skriver från terminalprompten, visa  anvisad manualsida:</p>
<div class="screen"><pre class="contents "><span class="cmd command">man sshd_config</span>
</pre></div>
<p class="para">
            There are many directives in the <span class="app application">sshd</span> configuration
	    file controlling such things as communication settings, and authentication modes.
	    The following are examples of configuration directives that can be changed by
	    editing the <span class="file filename">/etc/ssh/sshd_config</span> file.
            </p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents">
                <p class="para">Innan du redigerar konfigurationsfilen bör du göra en kopia av originalfilen och skydda den från skrivning så att du har kvar originalinställningarna som en referens och att återanvända om det blir nödvändigt.</p>
                <p class="para">Kopiera filen <span class="file filename">/etc/ssh/sshd_config</span> och skrivskydda den med följande kommandon som du skriver från en terminalprompt:</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo cp /etc/ssh/sshd_config /etc/ssh/sshd_config.original</span>
<span class="cmd command">sudo chmod a-w /etc/ssh/sshd_config.original</span>
</pre></div>
	    </div></div></div></div>
<p class="para">Följande är exempel på konfigurationsinställningar du kanske vill ändra på:</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
               <p class="para">För att få OpenSSH att lyssna på TCP-porten 2222 istället för standardporten 22, ändra raden Port så att den ser ut såhär:</p>
               <p class="para">Port 2222</p>
               </li>
<li class="list itemizedlist">
            <p class="para">För att få <span class="app application">sshd</span> att tillåta publika, nyckelbaserade inloggningsmetoder, lägg till eller ändra följande rad:</p>
               <p class="para">PubkeyAuthentication yes</p>
            <p class="para">
            If the line is already present, then ensure it is not commented out.
            </p>
            </li>
<li class="list itemizedlist">
             <p class="para">För att få OpenSSH-servern att visa innehållet i <span class="file filename">/etc/issue.net</span> som en inloggnings-banner, lägg till eller ändra följande rad:</p>
               <p class="para">Banner /etc/issue.net</p>
               <p class="para">I filen <span class="file filename">/etc/ssh/sshd_config</span>.</p>
             </li>
</ul></div>
<p class="para">Efter att du ändrat i filen <span class="file filename">/etc/ssh/sshd_config</span>, måste du spara den och starta om serverprogrammet <span class="app application">sshd</span> för att verkställa ändringarna. Du gör det genom att skriva följande kommando från terminalprompten:</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo systemctl restart sshd.service</span>
</pre></div>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents">
                  <p class="para">
                  Many other configuration directives for <span class="app application">sshd</span> are
	          available to change the server application's behavior to fit your needs.
		  Be advised, however, if your only method of access to a server is
		  <span class="app application">ssh</span>, and you make a mistake in configuring
		  <span class="app application">sshd</span> via the
		  <span class="file filename">/etc/ssh/sshd_config</span> file, you may find you
                  are locked out of the server upon restarting it. Additionally, if an incorrect configuration directive is supplied,
        	  the <span class="app application">sshd</span> server may refuse to start, so be extra careful when editing this file on a
		  remote server.
                  </p>
                </div></div></div></div>
</div></div>
</div></div>
<div class="sect2 sect" id="openssh-keys"><div class="inner">
<div class="hgroup"><h2 class="title">SSH-nycklar</h2></div>
<div class="region"><div class="contents">
<p class="para">
     SSH <span class="em emphasis">keys</span> allow authentication between two hosts without the need of a password.  SSH key authentication
     uses two keys, a <span class="em emphasis">private</span> key and a <span class="em emphasis">public</span> key.
     </p>
<p class="para">För att skapa nycklarna, skriv från en terminalprompt:</p>
<div class="screen"><pre class="contents "><span class="cmd command">ssh-keygen -t rsa</span>
</pre></div>
<p class="para">
     This will generate the keys using the <span class="em emphasis">RSA Algorithm</span>.  During the process you
     will be prompted for a password.  Simply hit <span class="em emphasis">Enter</span> when prompted to create the key.
     </p>
<p class="para">
     By default the <span class="em emphasis">public</span> key is saved in the file <span class="file filename">~/.ssh/id_rsa.pub</span>, while
     <span class="file filename">~/.ssh/id_rsa</span> is the <span class="em emphasis">private</span> key.  Now copy the <span class="file filename">id_rsa.pub</span> file
     to the remote host and append it to <span class="file filename">~/.ssh/authorized_keys</span> by entering:
     </p>
<div class="screen"><pre class="contents "><span class="cmd command">ssh-copy-id username@remotehost</span>
</pre></div>
<p class="para">Avslutningsvis, dubbelkontrollera tillstånden i filen <span class="file filename">authorized_keys</span>, enbart den verifierade användaren skall ha läs och skrivrättigheter. Om rättigheterna är felaktiga ändra dem genom att:</p>
<div class="screen"><pre class="contents "><span class="cmd command">chmod 600 .ssh/authorized_keys</span>
</pre></div>
<p class="para">Du skall nu kunna använda SSH till värden utan att behöva ange ett lösenord.</p>
</div></div>
</div></div>
<div class="sect2 sect" id="openssh-references"><div class="inner">
<div class="hgroup"><h2 class="title">Referenser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
          <p class="para">
          <a href="https://help.ubuntu.com/community/SSH" class="ulink" title="https://help.ubuntu.com/community/SSH">Ubuntu Wiki SSH</a> page.
          </p>
        </li>
<li class="list itemizedlist">
          <p class="para">
          <a href="http://www.openssh.org/" class="ulink" title="http://www.openssh.org/">OpenSSH:s webbplats</a>
          </p>
        </li>
<li class="list itemizedlist">
          <p class="para">
          <a href="https://wiki.ubuntu.com/AdvancedOpenSSH" class="ulink" title="https://wiki.ubuntu.com/AdvancedOpenSSH">Wikisida för avancerad OpenSSH-användning</a>
          </p>
        </li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="remote-administration.html" title="Fjärradministration">Föregående</a><a class="nextlinks-next" href="puppet.html" title="Puppet">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
