<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Tangentbord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 23.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 23.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Tangentbord</span></h1></div>
<div class="region">
<div class="contents pagewide">
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Region &amp; språk</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="keyboard-layouts.html.sv" title="Använd alternativa tangentbordslayouter">Använd alternativa tangentbordslayouter</a><span class="desc"> — Lägg till tangentbordslayouter och växla mellan dem.</span>
</li></ul></div>
</div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Hjälpmedel</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="a11y-stickykeys.html.sv" title="Aktivera klistriga tangenter">Aktivera klistriga tangenter</a><span class="desc"> — Mata in snabbtangenter en tangent i taget i stället för att hålla ner alla tangenterna på en gång.</span>
</li>
<li class="links ">
<a href="a11y-bouncekeys.html.sv" title="Aktivera tangentstuds">Aktivera tangentstuds</a><span class="desc"> — Ignorera snabbt repeterade tangenttryckningar på samma tangent.</span>
</li>
<li class="links ">
<a href="a11y-slowkeys.html.sv" title="Aktivera tröga tangenter">Aktivera tröga tangenter</a><span class="desc"> — Aktivera en fördröjning mellan tangenttryckning till det att bokstaven syns på skärmen.</span>
</li>
<li class="links ">
<a href="keyboard-osk.html.sv" title="Använd ett skärmtangentbord">Använd ett skärmtangentbord</a><span class="desc"> — Använd ett skärmtangentbord för att mata in text genom att klicka på knappar med musen eller en pekskärm.</span>
</li>
<li class="links ">
<a href="keyboard-nav.html.sv" title="Tangentbordsnavigation">Tangentbordsnavigation</a><span class="desc"> — Använd program och skrivbordet utan en mus.</span>
</li>
<li class="links ">
<a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?">Vad är <span class="key"><kbd>Super</kbd></span>-knappen?</a><span class="desc"> — <span class="key"><kbd>Super</kbd></span>-tangenten öppnar översiktsvyn <span class="gui">Aktiviteter</span>. Du kan vanligtvis hitta den intill <span class="key"><kbd>Alt</kbd></span>-tangenten på ditt tangentbord.</span>
</li>
<li class="links ">
<a href="keyboard-key-menu.html.sv" title="Vad är Windows-tangenten?">Vad är <span class="key"><kbd>Windows</kbd></span>-tangenten?</a><span class="desc"> — Tangenten <span class="key"><kbd>Meny</kbd></span> startar en snabbvalsmeny med tangentbordet snarare än med ett högerklick.</span>
</li>
</ul></div>
</div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Övriga ämnen</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar">Användbara tangentbordsgenvägar</a><span class="desc"> — Ta sig runt på skrivbordet med hjälp av tangentbordet.</span>
</li>
<li class="links ">
<a href="keyboard-cursor-blink.html.sv" title="Få tangentbordsmarkören att blinka">Få tangentbordsmarkören att blinka</a><span class="desc"> — Få insättningspunkten att blinka och kontrollera hur snabbt den blinkar.</span>
</li>
<li class="links ">
<a href="keyboard-repeat-keys.html.sv" title="Hantera repeterade tangenttryckningar">Hantera repeterade tangenttryckningar</a><span class="desc"> — Få tangentbordet att inte repetera bokstäver när du håller ner en tangent, eller ändra fördröjningen och hastigheten på repeterande tangenter.</span>
</li>
<li class="links ">
<a href="numeric-keypad.html.sv" title="Numeriskt tangentbord">Numeriskt tangentbord</a><span class="desc"> — Aktivera numeriska tangentbordet som standard.</span>
</li>
<li class="links ">
<a href="keyboard-shortcuts-set.html.sv" title="Ställ in tangentbordsgenvägar">Ställ in tangentbordsgenvägar</a><span class="desc"> — Definiera eller ändra snabbtangenter i inställningarna för <span class="gui">Tangentbord</span>.</span>
</li>
</ul></div>
</div></div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — Få GNOME att arbeta för dig, från hårdvarukontroll till sekretessinställningar.</span>
</li>
<li class="links ">
<a href="hardware.html.sv" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a><span class="desc"> — Konfigurera hårdvara och diagnostisera problem, inklusive skrivare, skärmar, diskar med mera.</span>
</li>
</ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
