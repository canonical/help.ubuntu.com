<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Kernel Crash Dump</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="installation.html" title="Installation">Installation</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="advanced-installation.html" title="Avancerad installation">Föregående</a><a class="nextlinks-next" href="package-management.html" title="Pakethantering">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Kernel Crash Dump</h1></div>
<div class="region">
<div class="contents"></div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="kernel-crash-dump.html#kernel-dump-introduction" title="Inledning">Inledning</a></li>
<li class="links"><a class="xref" href="kernel-crash-dump.html#kernel-crash-dump-mechanisms" title="Kernel Crash Dump Mechanism">Kernel Crash Dump Mechanism</a></li>
<li class="links"><a class="xref" href="kernel-crash-dump.html#Installation" title="Installation">Installation</a></li>
<li class="links"><a class="xref" href="kernel-crash-dump.html#kernel-dump-configuration" title="Konfiguration">Konfiguration</a></li>
<li class="links"><a class="xref" href="kernel-crash-dump.html#verification" title="Bekräftelse">Bekräftelse</a></li>
<li class="links"><a class="xref" href="kernel-crash-dump.html#kdump-testing" title="Testing the Crash Dump Mechanism">Testing the Crash Dump Mechanism</a></li>
<li class="links"><a class="xref" href="kernel-crash-dump.html#kdump-resources" title="Resurser">Resurser</a></li>
</ul></div>
<div class="sect2 sect" id="kernel-dump-introduction"><div class="inner">
<div class="hgroup"><h2 class="title">Inledning</h2></div>
<div class="region"><div class="contents"><p class="para">
        A Kernel Crash Dump refers to a portion of the contents of volatile memory (RAM) that is copied to disk whenever
         the execution of the kernel is disrupted. The following events can cause a kernel disruption :
         <div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist"><p class="para">Kernel Panic</p></li>
<li class="list itemizedlist"><p class="para">Non Maskable Interrupts (NMI)</p></li>
<li class="list itemizedlist"><p class="para">Machine Check Exceptions (MCE)</p></li>
<li class="list itemizedlist"><p class="para">Hardware failure</p></li>
<li class="list itemizedlist"><p class="para">Manual intervention</p></li>
</ul></div>
	 For some of those events (panic, NMI) the kernel will react automatically and trigger the crash dump mechanism through <span class="em emphasis">kexec</span>. In other situations a manual intervention is required in order to capture the memory.
	 
	 Whenever one of the above events occurs, it is important to find out the root cause in order to prevent it from happening again.  The cause can be determined by inspecting the copied memory contents.
        </p></div></div>
</div></div>
<div class="sect2 sect" id="kernel-crash-dump-mechanisms"><div class="inner">
<div class="hgroup"><h2 class="title">Kernel Crash Dump Mechanism</h2></div>
<div class="region"><div class="contents"><p class="para">
	When a kernel panic occurs, the kernel relies on the <span class="em emphasis">kexec</span> mechanism to quickly reboot a new instance of the kernel in a pre-reserved section of memory that had been allocated when the system booted (see below). This permits the existing memory area to remain untouched in order to safely copy its contents to storage.
        </p></div></div>
</div></div>
<div class="sect2 sect" id="Installation"><div class="inner">
<div class="hgroup"><h2 class="title">Installation</h2></div>
<div class="region"><div class="contents">
<p class="para">
      The kernel crash dump utility is installed with the following command:
      </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt-get install linux-crashdump</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="kernel-dump-configuration"><div class="inner">
<div class="hgroup"><h2 class="title">Konfiguration</h2></div>
<div class="region"><div class="contents">
<p class="para">
      Edit <span class="file filename">/etc/default/kdump-tools</span> by including the following line:
<div class="code"><pre class="contents ">USE_KDUMP=1
</pre></div>
      </p>
<p class="para">
      A reboot is then needed.
      </p>
</div></div>
</div></div>
<div class="sect2 sect" id="verification"><div class="inner">
<div class="hgroup"><h2 class="title">Bekräftelse</h2></div>
<div class="region"><div class="contents">
<p class="para">
      To confirm that the kernel dump mechanism is enabled, there are a few things to verify. First, confirm that
      the <span class="em emphasis">crashkernel</span> boot parameter is present (note: The following line has been split
      into two to fit the format of this document:
      </p>
<div class="screen"><pre class="contents "><span class="cmd command">cat /proc/cmdline</span>
<span class="output computeroutput">
BOOT_IMAGE=/vmlinuz-3.2.0-17-server root=/dev/mapper/PreciseS-root ro
 crashkernel=384M-2G:64M,2G-:128M
</span>
</pre></div>
<p class="para">
        The <span class="em emphasis">crashkernel</span> parameter has the following syntax: 
        <div class="code"><pre class="contents ">crashkernel=&lt;range1&gt;:&lt;size1&gt;[,&lt;range2&gt;:&lt;size2&gt;,...][@offset]
    range=start-[end] 'start' is inclusive and 'end' is exclusive.
        </pre></div>
	</p>
<p class="para"> 
So for the crashkernel parameter found in <span class="file filename">/proc/cmdline</span> we would have :
<div class="code"><pre class="contents ">crashkernel=384M-2G:64M,2G-:128M
</pre></div>
	</p>
<p class="para">The above value means:</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist"><p class="para">if the RAM is smaller than 384M, then don't reserve anything
       (this is the "rescue" case)</p></li>
<li class="list itemizedlist"><p class="para">if the RAM size is between 386M and 2G (exclusive), then reserve 64M</p></li>
<li class="list itemizedlist"><p class="para">if the RAM size is larger than 2G, then reserve 128M</p></li>
</ul></div>
<p class="para">
      Second, verify that the kernel has reserved the requested memory area for the kdump kernel by doing:
      </p>
<div class="screen"><pre class="contents "><span class="cmd command">dmesg | grep -i crash</span>
<span class="output computeroutput">
...
[    0.000000] Reserving 64MB of memory at 800MB for crashkernel (System RAM: 1023MB)
</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="kdump-testing"><div class="inner">
<div class="hgroup"><h2 class="title">Testing the Crash Dump Mechanism</h2></div>
<div class="region"><div class="contents">
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents">
	<p class="para">
	Testing the Crash Dump Mechanism will cause <span class="em emphasis">a system reboot.</span> In certain situations, this can
	cause data loss if the system is under heavy load. If you want to test the mechanism, make sure that the system
	is idle or under very light load.
	</p>
      </div></div></div></div>
<p class="para">
	Verify that the <span class="em emphasis">SysRQ</span> mechanism is enabled by looking at the value of the
	<span class="file filename">/proc/sys/kernel/sysrq</span> kernel parameter : 
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">cat /proc/sys/kernel/sysrq</span>
</pre></div>
<p class="para">
      If a value of <span class="em emphasis">0</span> is returned the feature is disabled. Enable it with the following command :
      </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo sysctl -w kernel.sysrq=1</span>
</pre></div>
<p class="para">
      Once this is done, you must become root, as just using <span class="cmd command">sudo</span> will not be sufficient. As the <span class="em emphasis">root</span>
      user, you will have to issue the command <span class="cmd command">echo c &gt; /proc/sysrq-trigger</span>. If you are using a network connection,
      you will lose contact with the system. This is why it is better to do the test while being connected to the system console. This has the 
      advantage of making the kernel dump process visible.
      </p>
<p class="para">
      A typical test output should look like the following :
      </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo -s</span>
[sudo] password for ubuntu: 
# <span class="cmd command">echo c &gt; /proc/sysrq-trigger</span>
[   31.659002] SysRq : Trigger a crash
[   31.659749] BUG: unable to handle kernel NULL pointer dereference at           (null)
[   31.662668] IP: [&lt;ffffffff8139f166&gt;] sysrq_handle_crash+0x16/0x20
[   31.662668] PGD 3bfb9067 PUD 368a7067 PMD 0 
[   31.662668] Oops: 0002 [#1] SMP 
[   31.662668] CPU 1 
....
</pre></div>
<p class="para">
      The rest of the output is truncated, but you should see the system rebooting and somewhere in the log, you will see the following line :
      <div class="screen"><pre class="contents ">Begin: Saving vmcore from kernel crash ...</pre></div>
      Once completed, the system will reboot to its normal operational mode. You will then find Kernel Crash Dump file in the <span class="file filename">/var/crash</span> directory :
      </p>
<div class="screen"><pre class="contents "><span class="cmd command">ls /var/crash</span>
linux-image-3.0.0-12-server.0.crash
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="kdump-resources"><div class="inner">
<div class="hgroup"><h2 class="title">Resurser</h2></div>
<div class="region"><div class="contents">
<p class="para">
      Kernel Crash Dump is a vast topic that requires good knowledge of the linux kernel. You can find more information on the topic here :
      </p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
              <p class="para">
              <a href="http://www.kernel.org/doc/Documentation/kdump/kdump.txt" class="ulink" title="http://www.kernel.org/doc/Documentation/kdump/kdump.txt">Kdump kernel documentation</a>.
              </p>
            </li>
<li class="list itemizedlist">
              <p class="para">
              <a href="http://people.redhat.com/~anderson/" class="ulink" title="http://people.redhat.com/~anderson/">The crash tool</a>
              </p>
            </li>
<li class="list itemizedlist">
              <p class="para">
              <a href="http://www.dedoimedo.com/computers/crash-analyze.html" class="ulink" title="http://www.dedoimedo.com/computers/crash-analyze.html">Analyzing Linux Kernel Crash</a> (Based on Fedora, it still gives a good walkthrough of kernel dump analysis)
              </p>
            </li>
</ul></div>
</div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="advanced-installation.html" title="Avancerad installation">Föregående</a><a class="nextlinks-next" href="package-management.html" title="Pakethantering">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
