<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Välj ett säkert lösenord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="user-accounts.html" title="Användarkonton">Users</a> › <a class="trail" href="user-accounts.html#passwords" title="Lösenord">Lösenord</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Välj ett säkert lösenord</span></h1></div>
<div class="region">
<div class="contents">
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">
      Make your passwords easy enough for you to remember, but very difficult 
      for others (including computer programs) to guess.
    </p></div></div></div></div>
<p class="p">
    Choosing a good password will help to keep your computer safe. If your 
    password is easy to guess, someone may figure it out and gain access to your 
    personal information.
  </p>
<p class="p">
    People could even use computers to systematically try to guess your 
    password, so even one that would be difficult for a human to guess might be 
    extremely easy for a computer program to crack. Here are some tips for 
    choosing a good password:
  </p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list">
<p class="p">
        Use a mixture of upper-case and lower-case letters, numbers, symbols, 
        and spaces in the password. This makes it more difficult to guess. There 
        are more symbols to choose from, so more possible passwords would have 
        to be checked by someone when trying to guess yours.
      </p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">
          A good method for choosing a password is to take the first letter of 
          each word in a phrase that you can remember. The phrase could be the 
          name of a movie, a book, a song, or an album. For example, "Flatland: 
          A Romance of Many Dimensions" would become F:ARoMD or faromd or f: 
          aromd.
        </p></div></div></div></div>
</li>
<li class="list"><p class="p">
        Make your password as long as possible. The more characters it contains, 
        the longer it should take for a person or computer to guess it.
      </p></li>
<li class="list"><p class="p">
        Do not use any words that appear in a standard dictionary in any 
        language. Password crackers will try these first. The most common 
        password is "password" -- people can guess passwords like this very 
        quickly!
      </p></li>
<li class="list"><p class="p">
        Do not use any personal information, such as a date, license plate 
        number, or any family member's name.
      </p></li>
<li class="list"><p class="p">
        Do not use any nouns.
      </p></li>
<li class="list">
<p class="p">
        Choose a password that can be typed quickly, to reduce the chance of 
        someone being able to make out what you have typed if they happen to be 
        watching you.
      </p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">
          Never write your passwords down anywhere. They can be found!
        </p></div></div></div></div>
</li>
<li class="list"><p class="p">
        Use different passwords for different things.
      </p></li>
<li class="list">
<p class="p">
        Use different passwords for different accounts.
      </p>
<p class="p">
        If you use the same password for all of your accounts, anyone who 
        guesses it will be able to access all of your accounts immediately.
      </p>
<p class="p">
        It can be difficult to remember lots of passwords. Though not as secure 
        as using a different passwords for everything, it may be easier to use 
        the same one for things that don't matter (like websites), and different 
        ones for important things (like your online banking account and your 
        email).
      </p>
</li>
<li class="list"><p class="p">
        Change your passwords regularly.
      </p></li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="user-accounts.html#passwords" title="Lösenord">Lösenord</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="user-changepassword.html" title="Välj ditt lösenord">Välj ditt lösenord</a><span class="desc"> — Keep your account secure by changing your password often
    in your account settings.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
