<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Dela ditt skrivbord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="sharing.html" title="Dela">Dela</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Dela ditt skrivbord</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan låta andra se och styra ditt skrivbord från en annan dator med ett skrivbordsvisningsprogram. Anpassa <span class="app">Skrivbordsdelning</span> för att låta andra komma åt ditt skrivbord, och ange säkerhetsinställningarna.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">I <span class="gui">Snabbstartspanelen</span>, öppna <span class="app">Skrivbordsdelning</span>.</p></li>
<li class="steps"><p class="p">För att låta andra se ditt skrivbord, välj <span class="gui">Låt andra användare se ditt skrivbord</span>. Detta betyder att andra kommer kunna försöka ansluta till din dator och se vad som visas på din skärm.</p></li>
<li class="steps"><p class="p">Fär att låta andra interagera med ditt skrivbord, välj <span class="gui">Låt andra användare styra ditt skrivbord</span>. Detta kan låta den andra personen flytta på din mus, köra program, och bläddra bland filer på din dator, beroende på aktuella säkerhetsinställningar.</p></li>
</ol></div></div></div>
</div>
<div id="security" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Säkerhet</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Det är viktigt att du funderar på den fulla vidden av vad varje säkerhetsalternativ innebär innan du ändrar det.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Bekräfta åtkomst till din maskin</dt>
<dd class="terms">
<p class="p">Om du vill kunna välja om någon ska kunna komma åt ditt skrivbord, välj <span class="gui">Du måste bekräfta varje åtkomst till den här maskinen</span>. Om du inaktiverar det här alternativet kommer du inte bli tillfrågad om du vill att någon ska kunna ansluta till din dator.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Detta alternativ är aktiverat som standard.</p></div></div></div></div>
</dd>
<dt class="terms">Aktivera lösenord</dt>
<dd class="terms">
<p class="p">För att kräva att andra använder lösenord när de ansluter till ditt skrivbord, välj <span class="gui">Kräv att användaren använder detta lösenord</span>. Om du inte använder det här alternativet kommer vem som helst kunna försöka se ditt skrivbord.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Detta alternativ är inaktiverat som standard, men du bör aktivera det och ställa in ett säkert lösenord.</p></div></div></div></div>
</dd>
<dt class="terms">Tillåt åtkomst till ditt skrivbord över internet</dt>
<dd class="terms">
<p class="p">Om din router har stöd för UPnP Internet Gateway-enhetprotokoll och det är aktiverat kan du tillåta att andra, som inte finns i ditt lokala nätverk, kan se ditt skrivbord. För att tillåta detta, välj <span class="gui">Ställ automatiskt in UPnP-router till att öppna och vidarebefordra portar</span>. Du kan annars justera din router manuellt.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Det här alternativet är avstängt som standard.</p></div></div></div></div>
</dd>
</dl></div></div></div>
</div></div>
</div></div>
<div id="notification-icon" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Visa ikon i notisfältet</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att kunna koppla bort någon som ser ditt skrivbord behöver du aktivera det här alternativet. Om du väljer <span class="gui">Alltid</span> kommer ikonen visas vare sig någon ser på ditt skrivbord eller inte.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om det här alternativet är avaktiverat är det möjligt för någon att ansluta till ditt skrivbord utan din vetskap, beroende på säkerhetsinställningarna.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="sharing.html" title="Dela">Dela</a><span class="desc"> — <span class="link"><a href="sharing-desktop.html" title="Dela ditt skrivbord">Skrivbordsdelning</a></span>, <span class="link"><a href="files-share.html" title="Dela ut och överför filer">Dela filer</a></span>...</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
