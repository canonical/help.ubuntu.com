<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Förhandsgranskningsinställningar för filhanterare</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 23.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a> » <a class="trail" href="nautilus-prefs.html.sv" title="Inställningar för filhanterare">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Förhandsgranskningsinställningar för filhanterare</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Filhanteraren skapar miniatyrbilder för att förhandsgranska bild-, video- och textfiler. Att skapa miniatyrbilder kan ta lång tid för stora filer eller över nätverk, så du kan styra när förhandsgranskning görs. Klicka på menyknappen i fönstrets övre högra hörn, välj <span class="gui">Inställningar</span> och gå sedan till avsnittet <span class="gui">Prestanda</span>.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Visa miniatyrbilder</span></dt>
<dd class="terms"><p class="p">Som standard görs förhandsgranskningar för <span class="gui">Bara på denna dator</span>, de på din dator eller anslutna externa hårddiskar. Du kan ställa in denna funktion till <span class="gui">Alla filer</span> eller <span class="gui">Aldrig</span>. Filhanteraren kan <span class="link"><a href="nautilus-connect.html.sv" title="Bläddra genom filer på en server eller nätverksutdelning">bläddra bland filer på andra datorer</a></span> över ett lokalt nätverk eller internet. Om du ofta bläddrar bland filer över ett lokalt nätverk och nätverket har en hög bandbredd kan det vara lämpligt att sätta förhandsgranskningsalternativet till <span class="gui">Alla filer</span>.</p></dd>
<dt class="terms"><span class="gui">Räkna antalet filer i mappar</span></dt>
<dd class="terms">
<p class="p">Om du visar filstorlekar i <span class="link"><a href="nautilus-list.html.sv" title="Kolumninställningar för listvy i Filer">listvykolumner</a></span> eller <span class="link"><a href="nautilus-display.html.sv#icon-captions" title="Ikonrubriker">ikonrubriker</a></span>, kommer mappar att visas tillsammans med antalet filer och mappar de innehåller. Att räkna antal objekt i en mapp kan gå långsamt, speciellt för väldigt stora mappar, eller över ett nätverk.</p>
<p class="p">Du kan slå av eller på denna funktion, eller slå på den endast för filer på din dator och lokala externa enheter.</p>
</dd>
</dl></div></div></div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="nautilus-prefs.html.sv" title="Inställningar för filhanterare">Inställningar för filhanterare</a><span class="desc"> — Visa och ställ in inställningar för filhanteraren.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-preview.html.sv" title="Förhandsgranska filer och mappar">Förhandsgranska filer och mappar</a><span class="desc"> — Visa och dölj snabbt förhandsgranskningar av dokument, bilder, videor och mera.</span>
</li></ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
