<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Redigera mappbokmärken</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#faq" title="Tips och frågor">Tips och frågor</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Redigera mappbokmärken</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Dina bokmärken är listade i sidopanelen i filhanteraren.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Lägg till ett bokmärke:</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna mappen (eller platsen) som du vill bokmärka.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Bokmärken</span> i menyraden och välj <span class="gui">Bokmärke för den här platsen</span>.</p></li>
</ol></div>
</div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Ta bort ett bokmärke:</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="gui">Bokmärken</span> i menyraden och välj <span class="gui">Bokmärken...</span> från programmenyn.</p></li>
<li class="steps"><p class="p">I fönstret <span class="gui">Bokmärken</span>, markera bokmärket du vill ta bort och klicka på <span class="key"><kbd>-</kbd></span>-knappen.</p></li>
</ol></div>
</div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Byt namn på ett bokmärke:</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="gui">Filer</span> i den övre raden och välj <span class="gui">Bokmärken</span> från programmenyn.</p></li>
<li class="steps"><p class="p">I fönstret <span class="gui">Bokmärken</span>, markera bokmärket du vill döpa om.</p></li>
<li class="steps">
<p class="p">I textrutan <span class="gui">Namn</span>, skriv in det nya namnet för bokmärket.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Att byta namn på ett bokmärke byter inte namn på mappen. Om du har bokmärken till två olika mappar på två olika platser, men som vart och ett har samma namn kommer bokmärkena att ha samma namn och du kommer inte att kunna skilja på dem. I dessa fall är det användbart att ge ett bokmärke ett namn annat än namnet på mappen som det pekar på.</p></div></div></div></div>
</li>
</ol></div>
</div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html#faq" title="Tips och frågor">Tips och frågor</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
