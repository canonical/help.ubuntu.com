<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ta bort filer och mappar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 21.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#common-file-tasks" title="Vanliga åtgärder">Vanliga åtgärder</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Ta bort filer och mappar</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Om du inte vill ha en fil eller mapp längre kan du ta bort den. När du tar bort ett objekt flyttas det till <span class="gui">Papperskorg</span> där det lagras tills du tömmer papperskorgen. Du kan <span class="link"><a href="files-recover.html.sv" title="Återskapa en fil från Papperskorgen">återställa objekt</a></span> i <span class="gui">Papperskorg</span> till deras originalplats om du bestämmer dig för att du behöver dem, eller om de togs bort av misstag.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">För att skicka en fil till papperskorgen:</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Markera objektet du önskar att placera i papperskorgen genom att klicka på det en gång.</p></li>
<li class="steps"><p class="p">Tryck <span class="key"><kbd>Delete</kbd></span> på ditt tangentbord. Alternativt, dra objektet till <span class="gui">Papperskorg</span> i sidopanelen.</p></li>
</ol></div>
</div></div>
<p class="p">Denna fil kommer att flyttas till papperskorgen och du kommer att kunna välja alternativet att <span class="gui">Ångra</span> borttagningen. <span class="gui">Ångra</span>-knappen kommer att visas under ett par sekunder. Om du väljer att <span class="gui">Ångra</span> kommer filen att återställas till dess ursprungliga plats.</p>
<p class="p">För att ta bort filer permanent och frigöra diskutrymme på din dator måste du tömma papperskorgen. För att tömma papperskorgen, högerklicka på <span class="gui">Papperskorg</span> i sidopanelen och välj <span class="gui">Töm papperskorgen</span>.</p>
</div>
<section id="permanent"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Ta bort en fil permanent</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Du kan ta bort en fil direkt, utan att behöva skicka den till papperskorgen först.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">För att permanent ta bort en fil:</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Markera objektet som du vill ta bort.</p></li>
<li class="steps"><p class="p">Tryck håll tangenten <span class="key"><kbd>Skift</kbd></span> nertryckt och tryck sedan på tangenten <span class="key"><kbd>Delete</kbd></span> på ditt tangentbord.</p></li>
<li class="steps"><p class="p">Eftersom du inte kan ångra detta kommer du att bli tillfrågad att bekräfta att du vill ta bort filen eller mappen.</p></li>
</ol></div>
</div></div>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Borttagna filer på en <span class="link"><a href="files.html.sv#removable" title="Flyttbara enheter och externa diskar">flyttbar enhet</a></span> är kanske inte synliga för andra operativsystem så som Windows eller Mac OS. Filerna är fortfarande där och kommer att vara tillgängliga när enheten återansluts till din dator.</p></div></div></div>
</div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html.sv#common-file-tasks" title="Vanliga åtgärder">Vanliga åtgärder</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="nautilus-behavior.html.sv#trash" title="Papperskorg">Papperskorgsinställningar för filhanterare</a></li>
<li class="links ">
<a href="files-recover.html.sv" title="Återskapa en fil från Papperskorgen">Återskapa en fil från Papperskorgen</a><span class="desc"> — Borttagna filer skickas normalt till Papperskorgen, men kan återställas.</span>
</li>
</ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
