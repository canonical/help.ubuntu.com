<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Handbok för Ubuntu-skrivbordet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" class="media media-inline" alt="Ubuntus logotyp"></span></span> Handbok för Ubuntu-skrivbordet</span></h1></div>
<div class="title" style="margin-bottom: 1.5em; margin-left: 0.8em"><span>Ubuntu 24.10</span></div><div class="region"><div class="contents pagewide">
<div class="links topiclinks"><div class="inner"><div class="region"><div class="tiles">
<div class="tile2 "><a class="ex-gnome-top" href="gnome-on-ubuntu.html.sv" title="Om GNOME i Ubuntu"><span class="ex-gnome-top-banner"></span><span class="ex-gnome-top-text"><span class="ex-gnome-top-title">Om GNOME i Ubuntu</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-top-desc">En lista över märkbara modifieringar av GNOME-skrivbordet i Ubuntu.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-top" href="shell-introduction.html.sv" title="Visuell överblick över GNOME"><span class="ex-gnome-top-banner"></span><span class="ex-gnome-top-text"><span class="ex-gnome-top-title">Visuell överblick över GNOME</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-top-desc">En visuell överblick över ditt skrivbord, systemraden, och översiktsvyn <span class="gui">Aktiviteter</span>.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-top" href="shell-exit.html.sv" title="Logga ut, stäng av eller växla användare"><span class="ex-gnome-top-banner"></span><span class="ex-gnome-top-text"><span class="ex-gnome-top-title">Logga ut, stäng av eller växla användare</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-top-desc">Lär dig hur du lämnar ditt användarkonto genom att logga ut, växla användare, och så vidare.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-top" href="shell-apps-open.html.sv" title="Starta program"><span class="ex-gnome-top-banner"></span><span class="ex-gnome-top-text"><span class="ex-gnome-top-title">Starta program</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-top-desc">Starta program från översiktsvyn <span class="gui">Aktiviteter</span>.</span></span></a></div>
<div class="tile2"></div>
</div></div></div></div>
<div class="links topiclinks"><div class="inner"><div class="region"><div class="tiles">
<div class="tile2 "><a class="ex-gnome-tile" href="shell-overview.html.sv" title="Ditt skrivbord"><span class="ex-gnome-tiles-banner"><img src="figures/tile-home.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Ditt skrivbord</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Arbeta med program, fönster och arbetsytor. Se dina möten och saker som är viktiga i systemraden.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="net.html.sv" title="Nätverk, webb &amp; e-post"><span class="ex-gnome-tiles-banner"><img src="figures/tile-net.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Nätverk, webb &amp; e-post</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Anslut till trådlösa och trådbundna nätverk. Håll dig säker med en VPN. Skapa en trådlös surfzon.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="media.html.sv" title="Ljud och media"><span class="ex-gnome-tiles-banner"><img src="figures/tile-media.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Ljud och media</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Hantera dina ljudenheter, använd dina mediafiler, anslut till externa enheter med mera.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="files.html.sv" title="Filer, mappar och sökning"><span class="ex-gnome-tiles-banner"><img src="figures/tile-files.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Filer, mappar och sökning</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Sök och hantera dina filer, oavsett om det är på din dator, på internet eller i säkerhetskopior.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="addremove.html.sv" title="Installera &amp; ta bort mjukvara"><span class="ex-gnome-tiles-banner"><img src="figures/tile-software.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Installera &amp; ta bort mjukvara</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Lägg till och ta bort applikationer och annan programvara. Hantera extra programvaruförråd.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="prefs.html.sv" title="Inställningar för användare och system"><span class="ex-gnome-tiles-banner"><img src="figures/tile-settings.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Inställningar för användare och system</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Få GNOME att arbeta för dig, från hårdvarukontroll till sekretessinställningar.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="hardware.html.sv" title="Maskinvara och drivrutiner"><span class="ex-gnome-tiles-banner"><img src="figures/tile-hardware.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Maskinvara och drivrutiner</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Konfigurera hårdvara och diagnostisera problem, inklusive skrivare, skärmar, diskar med mera.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="a11y.html.sv" title="Hjälpmedel"><span class="ex-gnome-tiles-banner"><img src="figures/tile-a11y.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Hjälpmedel</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Använd hjälpmedelsteknologier för att hjälpa till med speciella behov vad gäller syn, hörsel och rörlighet.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="tips.html.sv" title="Tips och tricks"><span class="ex-gnome-tiles-banner"><img src="figures/tile-tips.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Tips och tricks</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Få ut det mesta ur GNOME med dessa praktiska tips.</span></span></a></div>
<div class="tile2 "><a class="ex-gnome-tile" href="more-help.html.sv" title="Få mer hjälp"><span class="ex-gnome-tiles-banner"><img src="figures/tile-help.svg" width="" height="128"></span><span class="ex-gnome-tiles-text"><span class="ex-gnome-tiles-title">Få mer hjälp</span><span class="linkdiv-dash"> — </span><span class="ex-gnome-tiles-desc">Få tips om hur du använder denna guide, och ta kontakt med gemenskapen för mer hjälp.</span></span></a></div>
<div class="tile2"></div>
</div></div></div></div>
</div></div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
