<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Anslut en extern skärm till din bärbara dator</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="prefs-display.html" title="Visning och skärm">Visning och skärm</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Anslut en extern skärm till din bärbara dator</span></h1></div>
<div class="region">
<div class="contents"></div>
<div id="unity-steps" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ställ in en extern skärm</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att använda en extern skärm med din bärbara dator, anslut skärmen till datorn. Om ditt system inte känner igen den direkt, eller om du vill justera inställningarna:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="em">Systemmenyn</span> <span class="media"><span class="media media-image"><img src="figures/system-devices-panel.svg" class="media media-inline" alt="Kugghjulsikon"></span></span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Öppna <span class="gui">Skärmar</span>.</p></li>
<li class="steps"><p class="p">Klicka på bilden av den skärm du vill aktivera eller avaktivera, och växla mellan <span class="gui">PÅ/AV</span>.</p></li>
<li class="steps">
<p class="p">Som standard visas Programstartaren bara på primärskärmen. För att ändra vilken skärm som är ”primär”, ändra skärmen i den utfällbara rutan <span class="gui">Placering för Programstartaren</span>. Du skulle också kunna dra Programstartaren i förhandsgranskningen till skärmen du vill använda som primärskärm.</p>
<p class="p">Om du vill att Programstartaren ska visas på alla skärmar, ändra <span class="gui">Placering för Programstartaren</span> till <span class="gui">Alla skärmar</span>.</p>
</li>
<li class="steps">
<p class="p">För att ändra en skärms ”position”, klicka på den och dra den dit du vill ha den.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du vill att båda skärmarna ska visa samma bild, kryssa för rutan <span class="gui">Spegla skärmar</span>.</p></div></div></div></div>
</li>
<li class="steps"><p class="p">När du är nöjd med inställningarna, klicka på <span class="gui">Verkställ</span> och sedan <span class="gui">Behåll inställningarna</span>.</p></li>
<li class="steps"><p class="p">För att stänga <span class="gui">Skärmar</span>, klicka på <span class="gui">X:et</span> i det övre hörnet.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="sticky-edges" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Klistriga kanter</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Ett typiskt problem med två skärmar är att det är lätt för muspekaren att ”glida över” till den andra skärmen utan avsikt. Unitys funktion <span class="gui">Klistriga kanter</span> hjälper mot det problemet genom att kräva att du använder lite mer kraft för att flytta muspekaren från en skärm till en annan.</p>
<p class="p">Du kan stänga av <span class="gui">Klistriga kanter</span> om du inte tycker om funktionen.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs-display.html" title="Visning och skärm">Visning och skärm</a><span class="desc"> — <span class="link"><a href="look-background.html" title="Byt skrivbordsbakgrund">Bakgrund</a></span>, <span class="link"><a href="look-resolution.html" title="Ändra storlek och rotation för skärmen">storlek och orientering</a></span>, <span class="link"><a href="display-dimscreen.html" title="Ställ in skärmens ljusstyrka">ljusstyrka</a></span>...</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
