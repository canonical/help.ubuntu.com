<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Inställningar för användare och system</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 25.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Inställningar för användare och system</span></h1></div>
<div class="region">
<div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="user-accounts.html.sv" title="Användarkonton"><span class="title">Användarkonton</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till och ta bort användarkonton. Ändra lösenord. Ställ in administratörsbehörigheter.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="clock.html.sv" title="Datum och tid"><span class="title">Datum och tid</span><span class="linkdiv-dash"> — </span><span class="desc">Använd klockor och tidszoner, och håll koll på möten.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="prefs-sharing.html.sv" title="Dela-inställningar"><span class="title">Dela-inställningar</span><span class="linkdiv-dash"> — </span><span class="desc">Dela din skärm, eller dela media och andra filer över ett lokalt nätverk eller Bluetooth.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color.html.sv" title="Färghantering"><span class="title">Färghantering</span><span class="linkdiv-dash"> — </span><span class="desc">Kalibrera färgprofiler för skärmar, skrivare och andra enheter.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="media.html.sv#sound" title="Grundläggande ljud"><span class="title">Ljud</span><span class="linkdiv-dash"> — </span><span class="desc">Justera volymen för olika program, och konfigurera olika högtalare och mikrofoner.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm"><span class="title">Mus, styrplatta &amp; pekskärm</span><span class="linkdiv-dash"> — </span><span class="desc">Justera beteendet hos pekdon så att de uppfyller dina personliga krav.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="accounts.html.sv" title="Nätkonton"><span class="title">Nätkonton</span><span class="linkdiv-dash"> — </span><span class="desc">Anslut till dina konton med olika nättjänster.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="about.html.sv" title="Om"><span class="title">Om</span><span class="linkdiv-dash"> — </span><span class="desc">Visa information om ditt system.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="prefs-language.html.sv" title="Region &amp; språk"><span class="title">Region &amp; språk</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in dina föredragna språk, regioner, format och tangentbordslayouter.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="privacy.html.sv" title="Sekretessinställningar"><span class="title">Sekretessinställningar</span><span class="linkdiv-dash"> — </span><span class="desc">Lås din skärm, ta bort tillfälliga filer, och styr åtkomst till enheter som kameror och mikrofoner.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="quick-settings.html.sv" title="Snabbinställningar"><span class="title">Snabbinställningar</span><span class="linkdiv-dash"> — </span><span class="desc">Växla snabbt olika inställningar och välj enheter.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power.html.sv" title="Ström och batteri"><span class="title">Ström och batteri</span><span class="linkdiv-dash"> — </span><span class="desc">Visa din batteristatus och ändra strömsparinställningar.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="keyboard.html.sv" title="Tangentbord"><span class="title">Tangentbord</span><span class="linkdiv-dash"> — </span><span class="desc">Välj internationella tangentbordslayouter och använd hjälpmedelsfunktioner för tangentbordet.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="startup-applications.html.sv" title="Uppstartsprogram"><span class="title">Uppstartsprogram</span><span class="linkdiv-dash"> — </span><span class="desc">Välj vilka program som skall startas när du loggar in.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="prefs-display.html.sv" title="Visning och skärm"><span class="title">Visning och skärm</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in din bakgrund, konfigurera skärmar och hantera färgtemperaturer.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="wacom.html.sv" title="Wacom-ritplatta"><span class="title">Wacom-ritplatta</span><span class="linkdiv-dash"> — </span><span class="desc">Konfigurera din Wacom-ritplatta, inklusive spårningsläget och vilken skärm den är mappad till.</span></a></div>
</div>
</div></div></div></div></div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
