<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Användbara tangentbordsgenvägar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 25.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="keyboard.html.sv" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 25.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="keyboard.html.sv" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 25.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html.sv" title="Ditt skrivbord">Skrivbord</a> › <a class="trail" href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 25.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="tips.html.sv" title="Tips och tricks">Tips och tricks</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Användbara tangentbordsgenvägar</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Denna sida tillhandahåller en översikt över kortkommandon som kan hjälpa dig att använda ditt skrivbord och program mer effektivt. Om du inte kan använda en mus eller ett pekdon alls, se <span class="link"><a href="keyboard-nav.html.sv" title="Tangentbordsnavigation">Tangentbordsnavigation</a></span> för vidare information om hur man navigerar i användargränssnittet enbart med tangentbordet.</p>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="true"></div>
<div class="inner">
<div class="title title-table"><h2><span class="title">Ta sig runt på skrivbordet</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">tangenten <span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span></p></td>
<td><p class="p">Växla mellan översiktsvyn <span class="gui">Aktiviteter</span> och skrivbordet. I översiktsvyn kan du börja skriva för att omedelbart söka bland dina program, kontakter och dokument.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F2</kbd></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p">Visa kommandofönstret (för att snabbt köra kommandon).</p>
<p class="p">Använd piltangenterna för att snabbt komma åt tidigare körda kommandon.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-windows-switching.html.sv" title="Växla mellan fönster">Växla snabbt mellan fönster</a></span>. Håll ner <span class="key"><kbd>Skift</kbd></span> för omvänd ordning.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>`</kbd></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p">Växla mellan fönster från samma program, eller från det markerade programmet efter <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span>.</p>
<p class="p">Detta kortkommando använder <span class="key"><kbd>`</kbd></span> på amerikanska tangentbord, där tangenten <span class="key"><kbd>`</kbd></span> sitter ovanför <span class="key"><kbd>Tabb</kbd></span>. På alla andra tangentbord är kortkommandot <span class="key"><kbd>Super</kbd></span> samt tangenten ovanför <span class="key"><kbd>Tabb</kbd></span>.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Esc</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Växla mellan fönster i aktuell arbetsyta. Håll ner <span class="key"><kbd>Skift</kbd></span> för omvänd ordning.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Ge systemraden tangentbordsfokus. I översiktsvyn <span class="gui">Aktiviteter</span>, växla tangentbordsfokus mellan systemraden, snabbstartspanelen, fönsteröversiktsvyn, programlistan och sökfältet. Använd piltangenterna för att navigera.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>A</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Visa listan över program.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;">
<p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Up</kbd></span></span></p>
<p class="p">och</p>
<p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Down</kbd></span></span></p>
</td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-workspaces-switch.html.sv" title="Växla mellan arbetsytor">Växla mellan arbetsytor</a></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;">
<p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Up</kbd></span></span></p>
<p class="p">och</p>
<p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Down</kbd></span></span></p>
</td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-workspaces-movewindow.html.sv" title="Flytta ett fönster till en annan arbetsyta">Flytta det aktuella fönstret till en annan arbetsyta</a></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>←</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Flytta aktuellt fönster en skärm åt vänster.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>→</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Flytta aktuellt fönster en skärm åt höger.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Delete</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-exit.html.sv" title="Logga ut, stäng av eller växla användare">Visa dialogrutan Stäng av</a></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>L</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-exit.html.sv#lock-screen" title="Lås skärmen">Lås skärmen.</a></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>V</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Visa <span class="link"><a href="shell-notifications.html.sv#notificationlist" title="Aviseringslistan">aviseringslistan</a></span>. Tryck på <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>V</kbd></span></span> igen eller <span class="key"><kbd>Esc</kbd></span> för att stänga.</p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h2><span class="title">Vanliga redigeringsgenvägar</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>A</kbd></span></span></p></td>
<td><p class="p">Markera all text eller alla objekt i en lista.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>X</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Klipp ut markerad text eller objekt och placera dem i urklipp.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>C</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Kopiera markerad text eller objekt till urklipp.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>V</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Klistra in innehållet i urklipp.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Z</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Ångra senaste åtgärden.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>C</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Kopiera den markerade texten eller kommandona till urklipp i terminalen.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>V</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Klistra in innehållet i urklipp i terminalen.</p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h2><span class="title">Fånga från skärmen</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="key"><kbd>Print</kbd></span></p></td>
<td><p class="p"><span class="link"><a href="screen-shot-record.html.sv#screenshot" title="Ta en skärmbild">Starta skärmbildsverktyget.</a></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="screen-shot-record.html.sv#screenshot" title="Ta en skärmbild">Ta en skärmbild av ett fönster.</a></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="screen-shot-record.html.sv#screenshot" title="Ta en skärmbild">Ta en skärmbild av hela skärmen</a></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>R</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="screen-shot-record.html.sv#screencast" title="Gör en skärminspelning">Starta och stoppa en skärminspelning.</a></span></p></td>
</tr>
</table></div>
</div>
</div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a></li>
<li class="links ">
<a href="keyboard.html.sv" title="Tangentbord">Tangentbord</a><span class="desc"> — Välj internationella tangentbordslayouter och använd hjälpmedelsfunktioner för tangentbordet.</span>
</li>
<li class="links ">
<a href="tips.html.sv" title="Tips och tricks">Tips och tricks</a><span class="desc"> — Få ut det mesta ur GNOME med dessa praktiska tips.</span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="keyboard-shortcuts-set.html.sv" title="Ställ in tangentbordsgenvägar">Ställ in tangentbordsgenvägar</a><span class="desc"> — Definiera eller ändra snabbtangenter i inställningarna för <span class="gui">Tangentbord</span>.</span>
</li>
<li class="links ">
<a href="keyboard-nav.html.sv" title="Tangentbordsnavigation">Tangentbordsnavigation</a><span class="desc"> — Använd program och skrivbordet utan en mus.</span>
</li>
<li class="links ">
<a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?">Vad är <span class="key"><kbd>Super</kbd></span>-knappen?</a><span class="desc"> — <span class="key"><kbd>Super</kbd></span>-tangenten öppnar översiktsvyn <span class="gui">Aktiviteter</span>. Du kan vanligtvis hitta den intill <span class="key"><kbd>Alt</kbd></span>-tangenten på ditt tangentbord.</span>
</li>
<li class="links ">
<a href="keyboard-key-menu.html.sv" title="Vad är Windows-tangenten?">Vad är <span class="key"><kbd>Windows</kbd></span>-tangenten?</a><span class="desc"> — Tangenten <span class="key"><kbd>Meny</kbd></span> startar en snabbvalsmeny med tangentbordet snarare än med ett högerklick.</span>
</li>
</ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
