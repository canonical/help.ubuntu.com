<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Rapportera ett problem i Ubuntu</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 21.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="more-help.html.sv" title="Få mer hjälp">Få mer hjälp</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Rapportera ett problem i Ubuntu</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Om du hittar ett problem i Ubuntu kan du skicka in en <span class="em">felrapport</span>.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps">
<p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F2</kbd></span></span> och skriv <span class="input">ubuntu-bug namn-på-program</span></p>
<p class="p">Om du har ett hårdvaruproblem och inte vet vad det påverkade programmet heter, skriv bara <span class="input">ubuntu-bug</span></p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Om det av något skäl inte fungerar att använda <span class="cmd">ubuntu-bug</span>, <span class="link"><a href="https://help.ubuntu.com/community/ReportingBugs#Filing_bugs_manually_at_Launchpad.net" title="https://help.ubuntu.com/community/ReportingBugs#Filing_bugs_manually_at_Launchpad.net"> skicka in en felrapport manuellt</a></span> och hoppa till steg 4 i den här instruktionen.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Efter att du kör ett av ovanstående kommandon kommer Ubuntu samla in information om felet. Detta kan ta en stund. Granska den insamlade informationen om du vill. Klicka på <span class="gui">Skicka</span> för att fortsätta.</p></li>
<li class="steps"><p class="p">En ny flik kommer öppnas i webbläsaren för att fortsätta arbeta med felet. Ubuntu använder webbsidan <span class="app">Launchpad</span> för att hantera sina felrapporter. Om du inte har ett Launchpad-konto kommer du först behöva registrera ett för att skicka in din felrapport och få e-postuppdateringar om ärendet. Du kan göra det här genom att klicka på <span class="gui">Skapa nytt konto</span>.</p></li>
<li class="steps"><p class="p">Efter att du loggar in på Launchpad, beskriv problemet i sammanfattningsfältet.</p></li>
<li class="steps"><p class="p">Efter att du klickat på <span class="gui">Nästa</span> kommer Launchpad söka efter liknande felrapporter, för den händelse att felet du rapporterar redan har skickats in. Om felet redan har rapporterats kan du markera att det här felet påverkar dig också. Du kan också prenumerera på felrapporten för att ta emot uppdateringar om hur det går. Om felet inte redan har rapporterats, klicka på <span class="gui">Nej, jag behöver rapportera ett nytt fel</span>.</p></li>
<li class="steps">
<p class="p">Fyll i beskrivningsfältet med så mycket information du kan ge. Det är viktigt att du anger tre saker:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">Vad du förväntade dig skulle hända</p></li>
<li class="list"><p class="p">Vad som faktiskt hände</p></li>
<li class="list"><p class="p">Om möjligt, en minimal genomgång av de steg som ledde fram till felet, för steg 1 är "starta programmet"</p></li>
</ul></div></div></div>
</li>
<li class="steps"><p class="p">Din rapport kommer få ett ID-nummer, och dess tillstånd kommer uppdateras allt eftersom arbetet pågår. Tack för att du hjälper till att förbättra Ubuntu!</p></li>
</ol></div></div></div>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Om du för felmeddelandet "Det här är inte ett äkta Ubuntu-paket" innebär det att programmet du försöker felanmäla inte kommer från de officiella Ubuntu-arkiven. I så fall kan du inte använda Ubuntus inbyggda felrapporteringsverktyg.</p></div></div></div>
</div>
<p class="p">För mer information om hur du rapporterar fel i Ubuntu, läs den utförliga <span class="link"><a href="https://help.ubuntu.com/community/ReportingBugs" title="https://help.ubuntu.com/community/ReportingBugs">online-hjälpen</a></span>.</p>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="more-help.html.sv" title="Få mer hjälp">Få mer hjälp</a><span class="desc"> — <span class="link"><a href="about-this-guide.html.sv" title="Om denna handbok">Användningstips</a></span>, <span class="link"><a href="community-support.html.sv" title="Gemenskapssupport">få hjälp från gemenskapen</a></span>, <span class="link"><a href="get-involved.html.sv" title="Medverka till att förbättra den här handboken">hjälp till att förbättra handboken</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="get-involved.html.sv" title="Medverka till att förbättra den här handboken">Medverka till att förbättra den här handboken</a><span class="desc"> — Hur och var du ska rapportera problem med dessa hjälptexter.</span>
</li></ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
