<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Byobu</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="other-useful-applications.html" title="Ytterligare användbara program">Ytterligare användbara program</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="etckeeper.html" title="etckeeper">Föregående</a><a class="nextlinks-next" href="serverguide-appendix.html" title="Appendix">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Byobu</h1></div>
<div class="region">
<div class="contents">
<p class="para">
	    One of the most useful applications for any system administrator is an xterm multiplexor such as <span class="app application">screen</span> or
	    <span class="app application">tmux</span>.  It allows for the execution of multiple shells in one terminal. To make some of the advanced multiplexor
	    features more user-friendly and provide some useful information about the system, the <span class="app application">byobu</span> package was created.
	    It acts as a wrapper to these programs.  By default Byobu uses tmux (if installed) but this can be changed by the user.  
    </p>
<p class="para">
	    Invoke it simply with:
    </p>
<div class="screen"><pre class="contents "><span class="cmd command">byobu</span>
</pre></div>
<p class="para">
	Now bring up the configuration menu.  By default this is done by pressing the <span class="em emphasis">F9</span> key.  This will allow you to:
    </p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist"><p class="para">Visa hjälpmenyn</p></li>
<li class="list itemizedlist"><p class="para">Ändra Byobus bakgrundsfärg</p></li>
<li class="list itemizedlist"><p class="para">Ändra Byobus förgrundsfärg</p></li>
<li class="list itemizedlist"><p class="para">Växla statusnotifieringar</p></li>
<li class="list itemizedlist"><p class="para">Ändra tangentbordsgenvägar</p></li>
<li class="list itemizedlist"><p class="para">Ändra escape-sekvens</p></li>
<li class="list itemizedlist"><p class="para">Skapa nya fönster</p></li>
<li class="list itemizedlist"><p class="para">Hantera standardfönstren</p></li>
<li class="list itemizedlist"><p class="para">Byobu startas inte vid inloggning (aktivera)</p></li>
</ul></div>
<p class="para">
    The <span class="em emphasis">key bindings</span> determine such things as the escape sequence, new window, change window, etc.  There 
    are two key binding sets to choose from <span class="em emphasis">f-keys</span> and <span class="em emphasis">screen-escape-keys</span>.  If you wish to use the 
    original key bindings choose the <span class="em emphasis">none</span> set.
    </p>
<p class="para">
    <span class="app application">byobu</span> provides a menu which displays the Ubuntu release, processor information,
    memory information, and the time and date. The effect is similar to a desktop menu. 
    </p>
<p class="para">
    Using the <span class="em emphasis">"Byobu currently does not launch at login (toggle on)"</span> option will cause <span class="app application">byobu</span>
    to be executed any time a terminal is opened.  Changes made to <span class="app application">byobu</span> are on a per user basis, and will not 
    affect other users on the system.
    </p>
<p class="para">
    One difference when using byobu is the <span class="em emphasis">scrollback</span> mode.  Press the 
    <span class="em emphasis">F7</span> key to enter scrollback mode.  Scrollback mode allows you to navigate 
    past output using <span class="em emphasis">vi</span> like commands.  Here is a quick list of movement commands:
    </p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist"><p class="para"><span class="em emphasis">h</span> - Flytta markören ett tecken åt vänster</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">j</span> - Flytta markören ner en rad</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">k</span> - Flytta markören upp en rad</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">l</span> - Flytta markören ett tecken åt höger</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">0</span> - Flytta till början av nuvarande rad</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">$</span> - Flytta till slutet av nuvarande rad</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">G</span> - Flytta till den specificerade raden (standard till slutet av bufferten)</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">/</span> - Sök framåt</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">?</span> - Sök bakåt:</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">n</span> - Moves to the next match, either forward or backward</p></li>
</ul></div>
</div>
<div class="links sectionlinks" role="navigation"><ul><li class="links"><a class="xref" href="byobu.html#byobu-resources" title="Resurser">Resurser</a></li></ul></div>
<div class="sect2 sect" id="byobu-resources"><div class="inner">
<div class="hgroup"><h2 class="title">Resurser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
        <p class="para">För mer information om <span class="app application">screen</span> se webbplatsen för <a href="http://www.gnu.org/software/screen/" class="ulink" title="http://www.gnu.org/software/screen/">screen</a>.</p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        And the <a href="https://help.ubuntu.com/community/Screen" class="ulink" title="https://help.ubuntu.com/community/Screen">Ubuntu Wiki screen</a> page.
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        Also, see the <span class="app application">byobu</span> <a href="https://launchpad.net/byobu" class="ulink" title="https://launchpad.net/byobu">project page</a> for more
        information.
        </p>
      </li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="etckeeper.html" title="etckeeper">Föregående</a><a class="nextlinks-next" href="serverguide-appendix.html" title="Appendix">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
