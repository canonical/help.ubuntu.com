<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ansluta till nätet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="getting-started.html.sv" title="Komma igång">Börja med GNOME</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="gs-use-system-search.html.sv" title="Använd systemsökning">Föregående</a><a class="nextlinks-next" href="gs-browse-web.html.sv" title="Surfa på nätet">Nästa</a>
</div>
<div class="hgroup"><h1 class="title"><span class="title">Ansluta till nätet</span></h1></div>
<div class="region">
<div class="contents"><div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan se statusen för din nätverksuppkoppling på högersidan av systemraden.</p></div></div></div></div></div>
<div id="going-online-wired" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ansluta till ett trådbundet nätverk</span></h2></div>
<div class="region"><div class="contents">
<div class="media media-image"><div class="inner"><img src="gs-go-online1.svg" width="100%" class="media media-block" alt=""></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps">
<p class="p">Nätverksikonen på högersidan av systemraden visar att du är nedkopplad.</p>
<p class="p">Att vara nedkopplad kan ha flera orsaker: till exempel en nätverkskabel har kopplats ur, datorn har blivit inställd att köras i <span class="em">flygplansläge</span>, eller så finns det inga tillgängliga trådlösa nätverk i ditt närområde.</p>
<p class="p">Om du vill använda en trådbunden uppkoppling, koppla bara in en nätverkskabel för att ansluta till nätet. Datorn kommer att försöka ställa in nätverksuppkopplingen åt dig automatiskt.</p>
<p class="p">Medan datorn ställer in nätverksuppkopplingen åt dig så visar nätverksuppkopplingsikonen tre punkter.</p>
</li>
<li class="steps"><p class="p">När nätverksuppkopplingen har ställts in korrekt så ändras nätverksuppkopplingsikonen till symbolen för en nätverksansluten dator.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="going-online-wifi" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ansluta till ett trådlöst nätverk</span></h2></div>
<div class="region"><div class="contents">
<div class="media media-image"><div class="inner"><img src="gs-go-online2.svg" width="100%" class="media media-block" alt=""></div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">För att ansluta till ett trådlöst nätverk:</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="gui"><a href="shell-introduction.html.sv#yourname" title="Du och din dator">systemmenyn</a></span> på höger sida av systemraden.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Trådlöst nätverk ej anslutet</span>. Då kommer avdelningen om trådlösa nätverk att expanderas.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Välj nätverk</span>.</p></li>
</ol></div>
</div></div>
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan bara ansluta till ett trådlöst nätverk om din datorhårdvara har stöd för det och du befinner dig i ett område med täckning av minst ett trådlöst nätverk.</p></div></div></div></div>
<div class="media media-image"><div class="inner"><img src="gs-go-online3.svg" width="100%" class="media media-block" alt=""></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps" start="4"><li class="steps">
<p class="p">Från listan av tillgängliga trådlösa nätverk, välj det nätverk som du vill ansluta till och klicka <span class="gui">Koppla upp</span> för att bekräfta.</p>
<p class="p">Beroende på nätverkskonfigurationen, så kan du komma att bli ombedd att ange inloggningsuppgifter för nätverket.</p>
</li></ol></div></div></div>
</div></div>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="gs-use-system-search.html.sv" title="Använd systemsökning">Föregående</a><a class="nextlinks-next" href="gs-browse-web.html.sv" title="Surfa på nätet">Nästa</a>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="getting-started.html.sv" title="Komma igång">Börja med GNOME</a><span class="desc"> — Är GNOME nytt för dig? Lär dig hur du använder det.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a><span class="desc"> — <span class="link"><a href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlöst</a></span>, <span class="link"><a href="net-wired.html.sv" title="Trådbundna nätverk">trådbundet</a></span>, <span class="link"><a href="net-problem.html.sv" title="Nätverksproblem">anslutningsproblem</a></span>, <span class="link"><a href="net-browser.html.sv" title="Webbläsare">webbsurfning</a></span>, <span class="link"><a href="net-email.html.sv" title="E-post &amp; e-postprogramvara">e-postkonton</a></span>…</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
