<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="400" id="svg10075" version="1.1" ns1:version="0.48.4 r9939" ns2:docname="gs-web-browser1-firefox-classic.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,1.1342418,5.7016703,124.9606)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient5716-3-1">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-0-3"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-0-39"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient5716-3-1-9">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-0-3-4"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-0-39-8"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient5716-3-1-9-2">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-0-3-4-5"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-0-39-8-8"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-3-1" id="linearGradient31959" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-3-1-9" id="linearGradient31961" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-3-1-9-2" id="linearGradient31963" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-3-1-8-5-5" id="linearGradient5681-5" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient id="linearGradient5716-3-1-8-5-5">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-0-3-8-9-7"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-0-39-7-4-0"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient3962-1-1-9-5-4-2" id="radialGradient5559" gradientUnits="userSpaceOnUse" gradientTransform="matrix(0.66709696,0,0,0.66523581,301.76313,447.7745)" cx="18.247644" cy="15.716079" fx="18.247644" fy="15.716079" r="29.993349"/>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2">
      <ns0:stop id="stop3964-5-0-1-9-6-6" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient10586-8-2-5-1-6-0" id="linearGradient5561" gradientUnits="userSpaceOnUse" gradientTransform="matrix(0.12494518,0,0,0.125444,302.54321,448.90018)" x1="145.16281" y1="-41.407383" x2="144.42656" y2="46.077827"/>
    <ns0:linearGradient id="linearGradient10586-8-2-5-1-6-0" ns1:collect="always">
      <ns0:stop id="stop10588-8-7-5-8-3-4" offset="0" style="stop-color: rgb(172, 197, 237); stop-opacity: 1;"/>
      <ns0:stop id="stop10590-3-6-5-8-3-9" offset="1" style="stop-color: rgb(25, 59, 110); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5567" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:linearGradient id="linearGradient6868-5-7-5-4-3" ns1:collect="always">
      <ns0:stop id="stop6870-84-7-0-1-8" offset="0" style="stop-color: rgb(0, 0, 0); stop-opacity: 1;"/>
      <ns0:stop id="stop6872-0-5-0-7-1" offset="1" style="stop-color: rgb(0, 0, 0); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5565" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5563" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5573" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5571" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5569" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5579" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5577" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5575" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5585" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5583" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5581" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5591" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5589" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5587" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5597" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5595" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5593" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5603" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5601" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5599" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5609" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5607" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5605" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5615" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5613" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient5611" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient10599-4-0-8-1-6" id="radialGradient5617" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1.96261,0,0,1.09426,-74.6625,-21.1211)" cx="77.5625" cy="152.51079" fx="77.5625" fy="152.51079" r="13.03125"/>
    <ns0:linearGradient id="linearGradient10599-4-0-8-1-6" ns1:collect="always">
      <ns0:stop id="stop10601-9-3-6-7-5-5" offset="0" style="stop-color: rgb(255, 255, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop10603-3-0-1-5-1" offset="1" style="stop-color: rgb(255, 255, 255); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-3-1-8-5-5" id="linearGradient12974" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="677.05263" ns1:cy="217.78227" ns1:document-units="px" ns1:current-layer="layer2" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="2560" ns1:window-height="1408" ns1:window-x="2560" ns1:window-y="0" ns1:window-maximized="1" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-1092.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="830" x="-16" y="681.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-640)">
    <ns0:g id="g11020" transform="translate(-35,-52.36217)">
      <ns0:path transform="translate(2,453.36217)" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" ns2:ry="17" ns2:rx="17" ns2:cy="278" ns2:cx="120" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
      <ns0:text ns2:linespacing="125%" id="text11016" y="736.36218" x="122.29289" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan11018" ns2:role="line">1</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g id="g6333">
      <ns0:text ns2:linespacing="125%" id="text32728" y="742" x="84" style="font-size:12px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" xml:space="preserve"><ns0:tspan y="742" x="84" id="tspan32730" ns2:role="line">Program</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g transform="matrix(1.6306074,0,0,1.6324898,-290.27033,330.07988)" id="g3938">
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" id="rect3201" d="m 223.5,331.86218 0,-90 100,0" style="color:#000000;fill:#000000;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:1.83874416;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 224.5,261.36218 c 0,-2.48528 2.01471,-4.5 4.5,-4.5 l 109,0" style="fill:none;stroke:#000000;stroke-width:0.61291474px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" id="path3995"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 223.5,261.36218 c 0,-2.48528 2.01471,-4.5 4.5,-4.5 l 39,0" style="fill:none;stroke:#000000;stroke-width:1.83874416;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" id="path3995-8"/>
    </ns0:g>
    <ns0:g id="g5895" transform="matrix(1.3266261,0,0,1.2789155,-362.29125,797.60762)">
      <ns0:g transform="matrix(0.29958781,0,0,0.29170899,321.78845,-7.042621)" id="g5467">
        <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:7.7909255;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 464.46875,123.03125 0,0.125 c -0.44393,-0.0201 -0.89409,-0.0194 -1.3125,-0.0312 -0.0201,-5e-4 -0.0415,-6e-5 -0.0625,0 l 0,-0.0312 c -35.47303,0 -52.12084,18.17885 -58.53125,35.53125 -4.16563,11.27597 -2.56542,24.58143 -0.90625,38.0625 0.61719,5.01479 1.38934,10.3782 2.25,15.90625 0.0523,1.53427 0.0953,3.02176 0.0625,4.25 -0.48198,18.0321 -6.73844,40.14561 -6.375,53.75 0.67291,25.18859 14.15792,41.81557 32.09375,50.3125 0.28216,0.13367 0.55942,0.27661 0.84375,0.40625 20.53214,9.97483 44.84145,10.69846 64.53125,-2 17.00609,-9.04566 29.375,-25.39691 29.375,-48.71875 0,-13.60924 -5.89302,-35.7179 -6.375,-53.75 -0.19564,-7.31935 1.4375,-21.90625 1.4375,-21.90625 1.53635,-7.2428 2.64168,-15.026 2.34375,-22.59375 -0.004,-0.10339 0.005,-0.20919 0,-0.3125 -0.11179,-3.85613 -0.64084,-7.56265 -1.6875,-11.03125 -0.11795,-0.39089 -0.24268,-0.77221 -0.375,-1.15625 -0.10094,-0.32527 -0.172,-0.64602 -0.28125,-0.96875 -0.60655,-1.79171 -1.42373,-3.60933 -2.375,-5.40625 -0.0677,-0.13829 -0.15051,-0.26913 -0.21875,-0.40625 -11.84101,-23.79288 -32.00817,-30.03125 -54.4375,-30.03125 z" id="use3906-7-3"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="ccsccscsc" ns1:connector-curvature="0" id="path3896-9" d="m 471.25496,79.200587 5.30654,-28.587308 c 0.64849,-3.57802 1.26981,-7.661014 0.0259,-10.803791 -3.14471,-7.945086 -9.05873,-9.963605 -15.689,-9.963605 l -0.37971,0.0146 c -9.79602,0 -14.39338,5.126277 -16.16364,10.019502 l -3e-5,1e-6 c -1.15035,3.179726 -0.70845,6.93175 -0.25026,10.733293 0.74423,6.174786 2.22673,14.066104 3.59775,20.732961" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.38386175;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5509" d="m 460.5,28.862183 0,23" style="fill:none;stroke:#000000;stroke-width:0.38386175;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none"/>
      <ns0:rect ry="1.2794931" rx="1.1320361" y="35.253452" x="458.65408" height="11.488176" width="3.691813" id="rect5511" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:0.76772338;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 444,54.362183 c 5.14462,-1.307176 9.93443,-2.504355 16.4928,-2.499994 6.55838,-0.0044 11.34819,1.192829 16.49281,2.500005" style="fill:none;stroke:#000000;stroke-width:0.38386175;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" id="path5509-2-7"/>
    </ns0:g>
    <ns0:path style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0.95;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 207.77292,821.89434 -23.45593,-23.48299 8.0711,-8.08042 -29.97836,-2.3087 2.30604,30.01296 8.07109,-8.08041 39.95982,40.00596" id="rect12572" ns1:connector-curvature="0" ns2:nodetypes="ccccccc"/>
    <ns0:g transform="translate(343,-52.36217)" id="g31901">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path31903" ns2:cx="120" ns2:cy="278" ns2:rx="17" ns2:ry="17" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" transform="translate(2,453.36217)"/>
      <ns0:text xml:space="preserve" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="122.29289" y="736.36218" id="text31905" ns2:linespacing="125%"><ns0:tspan ns2:role="line" id="tspan31907" x="122.29289" y="736.36218">2</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g id="g5730-3" transform="matrix(1.3572719,0,0,1.3082544,494.71275,864.05898)">
      <ns0:g transform="matrix(0.29958781,0,0,0.29170899,381.78845,-7.042639)" id="g5467-6-5-7">
        <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:7.61561155;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 464.46875,123.03125 0,0.125 c -0.44393,-0.0201 -0.89409,-0.0194 -1.3125,-0.0312 -0.0201,-5e-4 -0.0415,-6e-5 -0.0625,0 l 0,-0.0312 c -35.47303,0 -52.12084,18.17885 -58.53125,35.53125 -4.16563,11.27597 -2.56542,24.58143 -0.90625,38.0625 0.61719,5.01479 1.38934,10.3782 2.25,15.90625 0.0523,1.53427 0.0953,3.02176 0.0625,4.25 -0.48198,18.0321 -6.73844,40.14561 -6.375,53.75 0.67291,25.18859 14.15792,41.81557 32.09375,50.3125 0.28216,0.13367 0.55942,0.27661 0.84375,0.40625 20.53214,9.97483 44.84145,10.69846 64.53125,-2 17.00609,-9.04566 29.375,-25.39691 29.375,-48.71875 0,-13.60924 -5.89302,-35.7179 -6.375,-53.75 -0.19564,-7.31935 1.4375,-21.90625 1.4375,-21.90625 1.53635,-7.2428 2.64168,-15.026 2.34375,-22.59375 -0.004,-0.10339 0.005,-0.20919 0,-0.3125 -0.11179,-3.85613 -0.64084,-7.56265 -1.6875,-11.03125 -0.11795,-0.39089 -0.24268,-0.77221 -0.375,-1.15625 -0.10094,-0.32527 -0.172,-0.64602 -0.28125,-0.96875 -0.60655,-1.79171 -1.42373,-3.60933 -2.375,-5.40625 -0.0677,-0.13829 -0.15051,-0.26913 -0.21875,-0.40625 -11.84101,-23.79288 -32.00817,-30.03125 -54.4375,-30.03125 z" id="use3906-7-3-7-4-1"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="ccsccscsc" ns1:connector-curvature="0" id="path3896-9-3-4-3" d="m 531.25496,79.200569 5.30654,-28.587308 c 0.64849,-3.57802 1.26981,-7.661014 0.0259,-10.803791 -3.14471,-7.945086 -9.05873,-9.963605 -15.689,-9.963605 l -0.37971,0.0146 c -9.79602,0 -14.39338,5.126277 -16.16364,10.019502 l -3e-5,10e-7 c -1.15035,3.179726 -0.70845,6.93175 -0.25026,10.733293 0.74423,6.174786 2.22673,14.066104 3.59775,20.732961" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.3752239;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path style="color:#000000;fill:#000000;stroke:none;stroke-width:3.00118113;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 520.5,28.874983 c -10.60524,0.01066 -15.58145,5.286996 -17.5,10.34375 -1.24797,3.289302 -0.77832,7.192451 -0.28125,11.125 0.15991,1.265137 0.37727,2.617453 0.59375,4 0.23237,0.0044 0.44738,0.03125 0.6875,0.03125 5.14462,-1.307176 9.93813,-2.504358 16.5,-2.5 l 0,-23 z" id="use3906-7-3-7-6-8-6-2" ns1:connector-curvature="0"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5509-5-9-7" d="m 520.5,28.862165 0,23" style="fill:none;stroke:#000000;stroke-width:0.3752239;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none"/>
      <ns0:rect ry="1.1118219" rx="1.1118219" y="35.241211" x="518.64331" height="11.488283" width="3.7133853" id="rect5511-0-2-1" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:0.75044769;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 503.99999,54.362165 c 5.14462,-1.307176 9.93443,-2.504355 16.4928,-2.499994 6.55838,-0.0044 11.34819,1.192829 16.49281,2.500005" style="fill:none;stroke:#000000;stroke-width:0.3752239;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" id="path5509-2-7-3-8-9"/>
    </ns0:g>
    <ns0:g transform="matrix(1.6699552,0,0,1.6699552,331.11105,831.90571)" id="g4614-7">
      <ns0:path style="fill:none;stroke:#000000;stroke-width:0.59834695;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 501.50039,55.861789 -4,0" id="path5939-2-0" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="21.49961"/>
      <ns0:path ns1:transform-center-y="-5.5645085" style="fill:none;stroke:#000000;stroke-width:0.59834695;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 502.16482,50.814919 -3.8637,-1.035277" id="path5939-2-4-6" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="20.76703"/>
      <ns0:path ns1:transform-center-y="-10.749805" style="fill:none;stroke:#000000;stroke-width:0.59834695;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 504.11284,46.112031 -3.4641,-2" id="path5939-2-4-0-2" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="18.61921"/>
      <ns0:path ns1:transform-center-y="-15.202521" style="fill:none;stroke:#000000;stroke-width:0.59834695;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="M 507.21169,42.073487 504.38327,39.24506" id="path5939-2-4-0-9-6" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="15.20252"/>
      <ns0:path ns1:transform-center-y="-18.61921" style="fill:none;stroke:#000000;stroke-width:0.59834695;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 511.25019,38.974664 -1.99999,-3.4641" id="path5939-2-4-0-9-1-7" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="10.749805"/>
      <ns0:path ns1:transform-center-y="-20.76703" style="fill:none;stroke:#000000;stroke-width:0.59834695;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 515.95313,37.026669 -1.03527,-3.8637" id="path5939-2-4-0-9-1-9-6" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="5.564505"/>
      <ns0:path ns1:transform-center-y="5.564509" style="fill:none;stroke:#000000;stroke-width:0.59834695;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 502.16482,60.908708 -3.8637,1.035274" id="path5939-2-4-4-7" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="20.76703"/>
    </ns0:g>
    <ns0:path style="color:#000000;fill:#000000;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 1071.1969,979.30312 0,-6.22187 m 0,-9.89844 0,-10.18125 m 0,-7.63594 0,-143.66875" id="rect3201-9-0" ns1:connector-curvature="0" ns2:nodetypes="cccccc"/>
    <ns0:path style="color:#000000;fill:none;stroke:#000000;stroke-width:0.99999988;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 1070.6313,937.72968 0,-128.11406 42.4218,0 c 3.1336,0 5.6563,2.52269 5.6563,5.65625 l 0,130.94219 m 0,6.7875 0,6.50469 m 0,3.67656 0,4.525" id="rect8340-2" ns1:connector-curvature="0" ns2:nodetypes="ccssccccc"/>
    <ns0:rect y="812.25208" x="1075.7146" height="39.608391" width="39.608391" id="rect8342-8-7-0" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.5;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" rx="2" ry="2"/>
    <ns0:path style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:1;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;fill-opacity:1" d="m 510.5,754.40625 -8.15625,8.15625 -12.8125,0 c -2.77,0 -5,2.23 -5,5 l 0,247 c 0,2.77 2.23,5 5,5 l 294,0 c 2.77,0 5,-2.23 5,-5 l 0,-247 c 0,-2.77 -2.23,-5 -5,-5 l -264.875,0 -8.15625,-8.15625 z" id="rect12158" ns1:connector-curvature="0"/>
    <ns0:g id="g5884-7" transform="matrix(1.13125,0,0,1.13125,239.7125,418.37778)">
      <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:2.65193367;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 340.78549,368.86218 -3.28539,3 -10e-4,26 23,0 -10e-4,-26 -3.28538,-3 -16.42693,0 z" id="rect2846-2-0-5" ns2:nodetypes="ccccccc"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccc" id="path4185-68-9-7-8" d="m 346.5,379.86218 0,1 5,0 0,-1" style="fill:none;stroke:#000000;stroke-width:0.88397789px;stroke-linecap:round;stroke-linejoin:round;stroke-opacity:1;display:inline;enable-background:new"/>
      <ns0:path ns2:nodetypes="ccccccc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-6-9" d="m 340.5,376.48718 0,-1.625 17,0 0,2.75 m 0,6.25 -17,0 0,-3.625" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.44198895;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cccccc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-3-4-8" d="m 357.5,385.86218 0,9 -17,0 m 0,-4.125 0,-4.875 11.6875,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.44198895;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccc" id="path4185-68-9-7-5-7" d="m 346.5,390.86218 0,1 5,0 0,-1" style="fill:none;stroke:#000000;stroke-width:0.88397789px;stroke-linecap:round;stroke-linejoin:round;stroke-opacity:1;display:inline;enable-background:new"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-6-4-5" d="m 340.5,372.86218 17,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.44198895;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:g>
    <ns0:g id="g5600-4" transform="matrix(1.13125,0,0,1.13125,239.7125,364.62778)">
      <ns0:path ns2:nodetypes="ccccccccccccc" id="rect2846-7-2-9-3-1-8-2" d="m 343.45832,368.86218 c -1.40839,0 -2.63187,0.7282 -3.2858,1.81251 l -1.08919,2.50961 c -0.37007,0.61442 -0.58333,1.32862 -0.58333,2.09134 l 0,18.40386 c 0,2.3172 1.95126,4.18268 4.37498,4.18268 l 12.25003,0 c 2.42373,0 4.37499,-1.86548 4.37499,-4.18268 l 0,-18.40386 c 0,-0.76272 -0.21325,-1.47692 -0.58333,-2.09134 l -1.08918,-2.50961 c -0.65395,-1.08431 -1.87742,-1.81251 -3.28582,-1.81251 l -11.08335,0 z" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:2.65193343;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#000000;stroke:#000000;stroke-width:0.44198892;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 349.00003,375.61218 c -1.46798,0 -2.80875,0.49981 -3.88406,1.33645 l -0.66823,0 c -0.25452,0 -0.45941,0.2049 -0.45941,0.45941 l 0,0.66823 c -0.83664,1.07531 -1.33645,2.41609 -1.33645,3.88406 0,1.46797 0.49981,2.80874 1.33645,3.88406 l 0,0.66822 c 0,0.25451 0.20489,0.45941 0.45941,0.45941 l 0.66823,0 c 1.07531,0.83663 2.41608,1.33645 3.88406,1.33645 1.46797,0 2.80874,-0.49982 3.88406,-1.33645 l 0.66821,0 c 0.25452,0 0.45942,-0.2049 0.45942,-0.45941 l 0,-0.66822 c 0.83664,-1.07532 1.33645,-2.41609 1.33645,-3.88406 0,-1.46797 -0.49981,-2.80875 -1.33645,-3.88406 l 0,-0.66823 c 0,-0.25451 -0.2049,-0.45941 -0.45942,-0.45941 l -0.66821,0 c -1.07532,-0.83664 -2.41609,-1.33645 -3.88406,-1.33645 z" id="path3861-6-2-2-7-4-1-1" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:0.88397789;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 349,376.96032 c -2.76142,0 -4.99998,2.23858 -4.99998,5 0,2.76142 2.23856,5 4.99998,5 2.76143,0 5,-2.23858 5,-5 0,-2.76142 -2.23857,-5 -5,-5 z" id="path3861-6-4-8-5-2-0-1" ns2:nodetypes="csssc" ns1:connector-curvature="0"/>
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path3861-6-1-6-2-1-0-0" ns2:cx="143.75" ns2:cy="155.25" ns2:rx="63.25" ns2:ry="63.25" d="m 207,155.25 c 0,34.93201 -28.31799,63.25 -63.25,63.25 C 108.81799,218.5 80.5,190.18201 80.5,155.25 80.5,120.31799 108.81799,92 143.75,92 178.68201,92 207,120.31799 207,155.25 z" transform="matrix(0.03324596,0,0,0.03324596,344.2209,376.79887)"/>
      <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path3861-6-1-3-8-2-2" ns2:cx="143.75" ns2:cy="155.25" ns2:rx="63.25" ns2:ry="63.25" d="m 207,155.25 c 0,34.93201 -28.31799,63.25 -63.25,63.25 C 108.81799,218.5 80.5,190.18201 80.5,155.25 80.5,120.31799 108.81799,92 143.75,92 178.68201,92 207,120.31799 207,155.25 z" transform="matrix(-0.02136966,0,0,-0.02078709,352.07189,385.03634)"/>
      <ns0:path ns2:nodetypes="csssc" ns1:connector-curvature="0" id="path5385-7-4-7-8-0" d="M 164.44918,225.50301 C 161.88194,223.3476 160.25,220.11438 160.25,216.5 c 0,-6.48935 5.26065,-11.75 11.75,-11.75 6.48935,0 11.75,5.26065 11.75,11.75 0,1.6575 -0.3432,3.23485 -0.96241,4.66485" style="color:#000000;fill:none;stroke:#000000;stroke-width:2.07734609;stroke-linecap:round;stroke-miterlimit:4;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(0.21276616,0,0,0.21276615,317.40422,346.29831)"/>
    </ns0:g>
    <ns0:g id="g8334" transform="matrix(1.13125,0,0,1.13125,689.4,478.31528)">
      <ns0:path ns2:nodetypes="cssssccc" ns1:connector-curvature="0" id="rect9426-5" d="m 344.5,436.42239 0,-13.13631 c 0,-0.78884 0.63171,-1.4239 1.4164,-1.4239 l 26.16723,0 c 0.78469,0 1.4164,0.63506 1.4164,1.4239 l 0,4.10735 m 0,1.96875 0,3" style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:2.65193367;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cccccccc" ns1:connector-curvature="0" id="rect9478-9" d="m 370.5,431.23718 0,2 m -22.99997,4.875 0,-3 m 0,-2 0,-7.25 22.99997,0 0,3.125" style="fill:none;stroke:#131616;stroke-width:0.44198895;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" id="path8330" d="m 349.5,427.86218 2.5,2 -2.5,2" style="fill:none;stroke:#000000;stroke-width:0.88397789px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path8332" d="m 353.58839,432.86218 3,0" style="fill:none;stroke:#000000;stroke-width:0.88397789px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1"/>
    </ns0:g>
    <ns0:g id="g30934" transform="matrix(0.55793991,0,0,0.55793991,337.25801,587.62468)">
      <ns0:path transform="matrix(0.96153846,0,0,0.96153846,133.63462,24.821622)" d="m 442.5,560.86218 c 0,16.2924 -13.2076,29.5 -29.5,29.5 -16.2924,0 -29.5,-13.2076 -29.5,-29.5 0,-16.2924 13.2076,-29.5 29.5,-29.5 16.2924,0 29.5,13.2076 29.5,29.5 z" ns2:ry="29.5" ns2:rx="29.5" ns2:cy="560.86218" ns2:cx="413" id="path30936" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6.24000025;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      <ns0:path style="fill:#ffffff;fill-opacity:1;stroke:none;display:inline" d="m 538.58035,543.84408 c -1.47456,-0.0645 -2.22819,0.0972 -2.21708,0.11066 0.0213,0.0285 6.13645,1.15986 7.20553,2.66049 0,0 -2.55107,0.0248 -5.09929,0.77601 -0.11531,0.0356 9.36682,1.17492 11.30712,10.8637 0,0 -1.0413,-2.284 -2.32796,-2.66051 0.84613,2.62977 0.5841,7.71838 -0.22171,10.19858 -0.10357,0.3189 -0.18623,-1.37501 -1.77366,-2.10625 0.5084,3.72199 -0.0214,9.57 -2.54966,11.19628 -0.19685,0.12664 1.55879,-5.84933 0.33242,-3.54732 -7.32057,11.46674 -15.98026,4.65062 -19.51035,2.21709 2.8333,0.7093 6.38645,0.24971 7.5381,-0.55428 1.75846,-1.2279 2.83489,-2.09673 3.76902,-1.88453 0.93373,0.21321 1.50118,-0.81354 0.776,-1.66279 -0.726,-0.85097 -2.49267,-1.96774 -4.8776,-1.33028 -1.68195,0.45006 -3.69122,1.9251 -6.87295,0 -2.71442,-1.64308 -2.37942,-2.48105 -2.37942,-3.33116 0,-0.85057 0.75869,-2.09674 2.10624,-1.88455 0.30187,0.0475 0.53472,0.0318 0.66512,0 0.65565,0.1497 1.26793,0.34196 1.88454,0.66512 0.0285,-0.79494 -0.10361,-3.0984 -0.55427,-4.36363 0.0376,0.0141 0.1025,0.0389 0.11065,0 0.13622,-0.62741 3.74164,-0.65222 4.87362,-2.11573 0.72381,-0.93514 0.49922,-2.82663 0.49922,-2.82663 l -3.54732,0 c -1.85719,0.008 -3.44958,-2.66355 -3.59881,-3.03896 0.40594,-2.22052 1.72443,-2.97804 3.59881,-4.05571 -1.41,-0.0107 -0.66942,0 -3.54736,0 -1.87562,0 -3.00521,1.28266 -3.59878,1.94947 -2.48519,-0.58837 -4.90045,-0.89487 -6.5998,-0.21603 -0.78485,-0.81378 -1.40488,-2.8398 -1.49655,-5.28064 0,0 -4.27402,2.62017 -3.82444,9.04969 -0.008,0.52869 -0.17701,0.75728 -0.2217,1.10855 -0.46333,0.81039 -0.55091,1.43637 -0.44341,1.33023 -0.23273,0.4834 -0.54596,1.00753 -0.776,1.66282 -0.0528,0.12841 -0.17557,0.16424 -0.22169,0.33239 -0.0318,0.11422 0.008,0.22631 0,0.3324 -0.40838,1.28055 -0.76324,3.48503 -1.10855,5.47216 0,0 0.44073,-1.82421 1.10855,-3.14424 -0.55478,1.92808 -0.9298,5.49744 -0.66512,9.68465 0,0 0.0533,-0.72468 0.22169,-1.77366 0.16495,2.84146 0.91966,6.12753 2.99306,9.75515 5.1845,9.07231 13.80792,13.08558 22.83596,12.30482 1.57912,-0.10501 3.17978,-0.38432 4.76672,-0.77601 21.03296,-5.195 18.73433,-31.14975 18.73433,-31.14975 l -0.55426,3.8799 c 0,0 -0.85656,-7.09386 -1.88451,-9.75515 -1.57545,-4.07792 -2.21254,-4.10751 -2.21709,-4.1016 1.05511,2.73945 0.77598,4.21244 0.77598,4.21244 0,0 -1.81902,-5.10598 -6.76209,-6.7621 -2.92707,-0.98019 -5.17669,-1.37661 -6.65125,-1.44109 z" id="path159-6-3" ns1:connector-curvature="0" ns2:nodetypes="sccccccccccsccccscccccscccccccccccccccccccccccccccs"/>
    </ns0:g>
    <ns0:g id="g12517-4-3" transform="matrix(1.4481746,0,0,1.4481746,-412.44396,377.66028)">
      <ns0:g style="stroke:#ffffff;stroke-width:3.45262241;stroke-miterlimit:4;stroke-dasharray:none" id="g12477-9-2-8" transform="translate(-3.6886788e-6,-1.0714912e-6)">
        <ns0:path ns1:transform-center-x="3.5" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-0-0-6" d="m 362.5,253.86218 -2,0" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none"/>
        <ns0:path ns1:transform-center-x="1.75" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-2-0-9" d="m 363.75,251.69712 -1,-1.73205" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:transform-center-y="-3.031085"/>
        <ns0:path ns1:transform-center-x="-1.75" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-7-1-0-1" d="m 366.25,251.69712 1,-1.73205" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:transform-center-y="-3.031085"/>
        <ns0:path ns1:transform-center-x="-3.5" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-7-0-2-0-0" d="m 367.5,253.86218 2,0" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none"/>
        <ns0:path ns1:transform-center-x="1.75" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-7-0-7-6-8-0" d="m 363.75,256.02724 -1,1.73205" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:transform-center-y="3.031085"/>
      </ns0:g>
      <ns0:g transform="translate(337.89511,250.27952)" ns1:label="#g5607" id="default-pointer-c-1-7-1-5" style="display:inline">
        <ns0:path style="color:#000000;fill:url(#linearGradient5681-5);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.69052446;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path5565-2-1-7-8" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path ns2:nodetypes="cccccccc" id="path6242-4-7-1-5" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.69052446;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:g id="g12477-99-7">
        <ns0:path ns1:transform-center-x="3.5" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-09-9" d="m 362.5,253.86218 -2,0" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none"/>
        <ns0:path ns1:transform-center-x="1.75" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-3-6" d="m 363.75,251.69712 -1,-1.73205" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:transform-center-y="-3.031085"/>
        <ns0:path ns1:transform-center-x="-1.75" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-7-4-9" d="m 366.25,251.69712 1,-1.73205" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:transform-center-y="-3.031085"/>
        <ns0:path ns1:transform-center-x="-3.5" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-7-0-73-6" d="m 367.5,253.86218 2,0" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none"/>
        <ns0:path ns1:transform-center-x="1.75" ns2:nodetypes="cc" ns1:connector-curvature="0" id="path5939-6-9-1-7-0-7-1-2" d="m 363.75,256.02724 -1,1.73205" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:transform-center-y="3.031085"/>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g12148" transform="matrix(1.6306074,0,0,1.6324898,105.72967,330.07988)">
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:1.83874416;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 223.5,331.86218 0,-90 100,0" id="path12150" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
      <ns0:path id="path12152" style="fill:none;stroke:#000000;stroke-width:0.61291474px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" d="m 224.5,261.36218 c 0,-2.48528 2.01471,-4.5 4.5,-4.5 l 109,0" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
      <ns0:path id="path12154" style="fill:none;stroke:#000000;stroke-width:1.83874416;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 223.5,261.36218 c 0,-2.48528 2.01471,-4.5 4.5,-4.5 l 39,0" ns1:connector-curvature="0" ns2:nodetypes="ccc"/>
    </ns0:g>
    <ns0:rect style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect12928" width="70" height="15" x="497" y="779" rx="0" ry="0"/>
    <ns0:rect ry="0" rx="0" y="799" x="497" height="15" width="78" id="rect12930" style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:rect style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect12932" width="56" height="15" x="497" y="819" rx="0" ry="0"/>
    <ns0:rect ry="0" rx="0" y="839" x="497" height="15" width="70" id="rect12934" style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:rect style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect12936" width="92" height="15" x="497" y="859" rx="0" ry="0"/>
    <ns0:rect ry="0" rx="0" y="879" x="497" height="15" width="70" id="rect12938" style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:rect style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect12940" width="95" height="15" x="497" y="982" rx="0" ry="0"/>
    <ns0:g transform="matrix(1.4481746,0,0,1.4481746,108.55604,542.66028)" id="g12942">
      <ns0:g transform="translate(-3.6886788e-6,-1.0714912e-6)" id="g12944" style="stroke:#ffffff;stroke-width:3.45262241;stroke-miterlimit:4;stroke-dasharray:none">
        <ns0:path style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 362.5,253.86218 -2,0" id="path12946" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="3.5"/>
        <ns0:path ns1:transform-center-y="-3.031085" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 363.75,251.69712 -1,-1.73205" id="path12948" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="1.75"/>
        <ns0:path ns1:transform-center-y="-3.031085" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 366.25,251.69712 1,-1.73205" id="path12950" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="-1.75"/>
        <ns0:path style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 367.5,253.86218 2,0" id="path12952" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="-3.5"/>
        <ns0:path ns1:transform-center-y="3.031085" style="fill:none;stroke:#ffffff;stroke-width:3.45262241;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 363.75,256.02724 -1,1.73205" id="path12954" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="1.75"/>
      </ns0:g>
      <ns0:g style="display:inline" id="g12956" ns1:label="#g5607" transform="translate(337.89511,250.27952)">
        <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccccccc" id="path12958" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" style="color:#000000;fill:url(#linearGradient12974);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.69052446;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate"/>
        <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.69052446;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path12960" ns2:nodetypes="cccccccc"/>
      </ns0:g>
      <ns0:g id="g12962">
        <ns0:path style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 362.5,253.86218 -2,0" id="path12964" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="3.5"/>
        <ns0:path ns1:transform-center-y="-3.031085" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 363.75,251.69712 -1,-1.73205" id="path12966" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="1.75"/>
        <ns0:path ns1:transform-center-y="-3.031085" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 366.25,251.69712 1,-1.73205" id="path12968" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="-1.75"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 367.5,253.86218 2,0" id="path12970" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="-3.5"/>
        <ns0:path ns1:transform-center-y="3.031085" style="fill:none;stroke:#000000;stroke-width:0.6899808;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 363.75,256.02724 -1,1.73205" id="path12972" ns1:connector-curvature="0" ns2:nodetypes="cc" ns1:transform-center-x="1.75"/>
      </ns0:g>
    </ns0:g>
    <ns0:rect ry="0" rx="0" y="893" x="663" height="15" width="76" id="rect13001" style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:rect style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect13003" width="50" height="15" x="663" y="843" rx="0" ry="0"/>
    <ns0:rect ry="0" rx="0" y="791" x="663" height="15" width="78" id="rect13005" style="color:#000000;fill:#babdb6;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:use x="0" y="0" ns4:href="#g6333" id="use6337" transform="translate(402,0)" width="840" height="400"/>
  </ns0:g>
</ns0:svg>
