<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använda programstartaren</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Använda programstartaren</span></h1></div>
<div class="region">
<div class="contents">
<div class="media media-image floatstart"><div class="inner"><img src="figures/unity-launcher-apps.png" class="media media-block" alt="Startarens ikoner"></div></div>
<p class="p"><span class="gui">Startaren</span> är en av de centrala komponenterna i skrivbordet Unity. När du loggar in på ditt skrivbord kommer den visas utmed skärmens vänstra sida. Startaren ger dig enkel åtkomst till program, arbetsytor, bärbara enheter, och papperskorgen.</p>
<p class="p">Om ett program som du vill börja använda finns på Programstartaren kan du klicka på programmets ikon, som då startas och är redo för att börja arbeta.</p>
<p class="p">För att läsa mer om Startaren, utforska någon av hjälprubrikerna om Startaren nedanför.</p>
</div>
<div id="launcher-using" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Använda Startaren</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="unity-launcher-menu.html" title="Startarens ikonmenyer"><span class="title">Startarens ikonmenyer</span><span class="linkdiv-dash"> — </span><span class="desc">Att högerklicka på en ikon på Programstartaren visar en meny med möjliga åtgärder.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-launcher-shapes.html" title="Vad betyder de olika formerna och färgerna på Startarens ikoner?"><span class="title">Vad betyder de olika formerna och färgerna på Startarens ikoner?</span><span class="linkdiv-dash"> — </span><span class="desc">Trianglarna visar dig vilka program som kör.</span></a></div>
</div></div></div></div></div>
</div></div>
<div id="launcher-customizing" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Anpassa Startaren</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-apps-favorites.html" title="Ändra vilka program som visas i Startaren"><span class="title">Ändra vilka program som visas i Startaren</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till, flytta, eller ta bort ofta använda programikoner på Startaren.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-launcher-change-autohide.html" title="Dölj Startaren automatiskt"><span class="title">Dölj Startaren automatiskt</span><span class="linkdiv-dash"> — </span><span class="desc">Visa <span class="gui">Startaren</span> bara när du behöver den.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="unity-launcher-change-size.html" title="Ändra storlek på ikonerna på Startaren"><span class="title">Ändra storlek på ikonerna på Startaren</span><span class="linkdiv-dash"> — </span><span class="desc">Gör ikonerna i Startaren större eller mindre.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
