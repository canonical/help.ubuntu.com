<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="500" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-go-online1.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns1:collect="always" id="linearGradient14901">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop14903"/>
      <ns0:stop style="stop-color:#000000;stop-opacity:0;" offset="1" id="stop14905"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2">
      <ns0:stop id="stop3964-5-0-1-9-6-6" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68893" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:linearGradient id="linearGradient6868-5-7-5-4-3" ns1:collect="always">
      <ns0:stop id="stop6870-84-7-0-1-8" offset="0" style="stop-color: rgb(0, 0, 0); stop-opacity: 1;"/>
      <ns0:stop id="stop6872-0-5-0-7-1" offset="1" style="stop-color: rgb(0, 0, 0); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68891" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68897" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68895" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68901" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68899" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68905" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68903" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68909" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68907" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68913" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68911" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68917" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68915" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68921" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68919" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68925" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68923" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath56767">
      <ns0:path ns2:nodetypes="ccccc" ns1:connector-curvature="0" id="path56769" d="m 228.45991,29.202459 833.57379,0 0,290.286071 c -330.23641,0 -408.68316,175.76954 -833.57379,175.76954 z" style="color:#000000;fill:#babdb6;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath14882">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:8.72566223;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path14884" ns2:cx="2246" ns2:cy="390" ns2:rx="482" ns2:ry="482" d="m 2728,390 a 482,482 0 1 1 -964,0 482,482 0 1 1 964,0 z" transform="matrix(0.35527386,0,0,0.35527386,119.03054,9.4159878)"/>
    </ns0:clipPath>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient14901" id="linearGradient14907" x1="532.43353" y1="187.53497" x2="532.43353" y2="314.62036" gradientUnits="userSpaceOnUse"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-2-7-1">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-4-6-6" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-1-4-3">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-5-5" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-3-9">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-5-4" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25942">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25944" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25946">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25948" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25950">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25952" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-9-6-0">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-1-6-2" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-6-4-2-8">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-19-7-4" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-8-2-8-7-5">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-9-2-7-6-1" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25960">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25962" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25964">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25966" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25968">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25970" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25972">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25974" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25976">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25978" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25980">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25982" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25984">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25986" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25988">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25990" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25992">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25994" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25996">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25998" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath26000">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect26002" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath26004">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect26006" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath24971-0" clipPathUnits="userSpaceOnUse">
      <ns0:rect y="-354.29291" x="624" height="93" width="276" id="rect24973-5" style="color:#000000;fill:none;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-2-7">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-4-6" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-1-4">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-5" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-3">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-5" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-1-7">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-9-9);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-5-6" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-5-5" id="radialGradient12116-6-2-9-3-0-9-9" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-5-5">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-4-1"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-8-15"/>
    </ns0:linearGradient>
    <ns0:clipPath id="clipPath4201-6-8-5-59">
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path4203-1-2-5-0" ns1:connector-curvature="0" d="m 101,177 0,5 2,0 0,2 1,0 0,-4 7,0 0,4 1,0 0,-2 2,0 0,-5 -13,0 z"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-9-6">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-1-6" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-6-4-2">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-19-7" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-8-2-8-7">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-9-2-7-6" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-3-7">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-75-13);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-6-5" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-7-2" id="radialGradient12116-6-2-9-3-0-75-13" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-7-2">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-8-92"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-04-00"/>
    </ns0:linearGradient>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-0-0">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-7-75);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-3-8" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-9-1" id="radialGradient12116-6-2-9-3-0-7-75" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-9-1">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-3-4"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-0-50"/>
    </ns0:linearGradient>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-4">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-3);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-0" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-77" id="radialGradient12116-6-2-9-3-0-3" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-77">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-87"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-7"/>
    </ns0:linearGradient>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath26963">
      <ns0:path style="color:#000000;fill:#204a87;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2.93785119;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 64,503 563,0 0,154 C 492.38459,818.58999 220.38142,629.28197 64,784 z" id="path26965" ns1:connector-curvature="0" ns2:nodetypes="ccccc"/>
    </ns0:clipPath>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient14901-1" id="linearGradient14907-7" x1="532.43353" y1="129.633" x2="532.43353" y2="177.87709" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient14901-1">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop14903-7"/>
      <ns0:stop style="stop-color:#000000;stop-opacity:0;" offset="1" id="stop14905-2"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(0.75098334,0,0,0.75098334,-170.84871,-42.430559)" y2="314.62036" x2="532.43353" y1="187.53497" x1="532.43353" gradientUnits="userSpaceOnUse" id="linearGradient27012" ns4:href="#linearGradient14901-1" ns1:collect="always"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-9">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9-8" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9-6" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6-7" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient14901" id="linearGradient27124" gradientUnits="userSpaceOnUse" x1="532.43353" y1="187.53497" x2="532.43353" y2="314.62036"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-7">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9-2" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4-5">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9-2" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2-8">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6-2" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient14901-1" id="linearGradient17826" gradientUnits="userSpaceOnUse" x1="532.43353" y1="129.633" x2="532.43353" y2="177.87709"/>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="300.20081" ns1:cy="205.65025" ns1:document-units="px" ns1:current-layer="layer2" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="2560" ns1:window-height="1401" ns1:window-x="2560" ns1:window-y="0" ns1:window-maximized="1" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="656" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-540)">
    <ns0:g id="g11020" transform="translate(-51,-143.36217)">
      <ns0:path transform="translate(2,453.36217)" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" ns2:ry="17" ns2:rx="17" ns2:cy="278" ns2:cx="120" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
      <ns0:text id="text11016" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan11018" ns2:role="line" style="font-size:14px;line-height:1.25">1</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g transform="matrix(0.49304709,0,0,0.49304709,-7.1085958,556.63869)" style="display:inline" id="g17515" ns1:export-filename="/home/jimmac/gfx/redhat/redhat-ux/Products/RHEL/RHEL7/video-jingles/tex/overview.png" ns1:export-xdpi="90" ns1:export-ydpi="90" clip-path="url(#clipPath56767)">
      <ns0:path ns2:nodetypes="ccccccc" ns1:connector-curvature="0" id="rect10989-4" d="m 239.06066,57.414214 800.87864,0 0,51.485276 c 0,0 -4.0279,-10.606597 -11.0989,-10.96015 L 249,99 c -4.59619,-0.353553 -9.93934,5.5 -9.93934,5.5 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:g transform="translate(11,0)" id="g10976-7">
        <ns0:path style="color:#000000;fill:none;stroke:url(#linearGradient27124);stroke-width:3;stroke-miterlimit:4;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 229,658 0,-600 800,0 0,67.36502" id="rect10923-0" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
        <ns0:path id="path10955-1" style="fill:none;stroke:#000000;stroke-width:2.37319922px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" d="m 1028.199,108.766 c 0,-5.89806 -4.7813,-10.6794 -10.6794,-10.6794 l -777.99931,0 c -5.89809,0 -10.6794,4.78134 -10.6794,10.6794" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
        <ns0:text id="text10968-2" y="86.187378" x="1014.3748" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="86.187378" x="1014.3748" id="tspan10970-0" ns2:role="line" style="font-size:21.26189423px;line-height:1.25">Maria Johansson</ns0:tspan></ns0:text>
        <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none" x="628.8465" y="86.187378" id="text10972-5"><ns0:tspan ns2:role="line" id="tspan10974-5" x="628.8465" y="86.187378" style="font-size:21.26189423px;line-height:1.25">14:30</ns0:tspan></ns0:text>
        <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="238.05931" y="86.187378" id="text56758"><ns0:tspan ns2:role="line" id="tspan56760" x="238.05931" y="86.187378" style="font-size:21.26189423px;line-height:1.25">Aktiviteter</ns0:tspan></ns0:text>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g14886" transform="matrix(0.72370712,0,0,0.72370712,-966.69401,132.94511)">
      <ns0:g transform="matrix(1.6234335,0,0,1.6234335,645.35105,529.77601)" style="display:inline" id="g14053" ns1:export-filename="/home/jimmac/gfx/redhat/redhat-ux/Products/RHEL/RHEL7/video-jingles/tex/overview.png" ns1:export-xdpi="90" ns1:export-ydpi="90" clip-path="url(#clipPath14882)">
        <ns0:path ns2:nodetypes="ccccccc" ns1:connector-curvature="0" id="path14055" d="m 239.06066,57.414214 800.87864,0 0,51.485276 c 0,0 -4.0279,-10.606597 -11.0989,-10.96015 L 249,99 c -4.59619,-0.353553 -9.93934,5.5 -9.93934,5.5 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:g transform="translate(11,0)" id="g14057">
          <ns0:rect style="color:#000000;fill:none;stroke:url(#linearGradient14907-7);stroke-width:1.38776851;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect14059" width="800" height="600" x="229" y="58.307991"/>
          <ns0:path id="path14061" style="fill:none;stroke:#000000;stroke-width:1.09781706px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" d="m 1028.815,108.766 c 0,-5.89806 -4.7813,-10.6794 -10.6794,-10.6794 l -777.99933,0 c -5.89809,0 -10.6794,4.78134 -10.6794,10.6794" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
        </ns0:g>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g27126" transform="translate(0,127.70887)">
      <ns0:g id="g15031" transform="translate(-51,24.637831)">
        <ns0:path transform="translate(2,453.36217)" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" ns2:ry="17" ns2:rx="17" ns2:cy="278" ns2:cx="120" id="path15033" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
        <ns0:text id="text15035" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan15037" ns2:role="line" style="font-size:14px;line-height:1.25">2</ns0:tspan></ns0:text>
      </ns0:g>
    </ns0:g>
    <ns0:rect style="color:#000000;fill:none;stroke:#000000;stroke-width:1.79821837;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:1.79821915, 1.79821915;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect27120" width="37.297157" height="37.297157" x="590.11682" y="590.58606" rx="5.4661207" ry="5.4661207"/>
    <ns0:g style="display:inline" ns1:label="audio-volume-medium" transform="matrix(1.333369,0,0,1.333369,604.00453,310.0695)" id="g5525">
      <ns0:path ns1:connector-curvature="0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none" d="m 20,222 h 2.484375 L 25.453129,219 26,219.0156 v 11 l -0.475297,8.3e-4 L 22.484375,227 H 20 Z" id="path5533" ns2:nodetypes="ccccccccc"/>
      <ns0:rect ns1:label="audio-volume-high" y="217" x="20" height="16" width="16" id="rect5535" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none"/>
      <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3718-5" style="display:inline;fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:type="arc" clip-path="url(#clipPath6279-7-9-7)"/>
      <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" ns2:type="arc" style="display:inline;fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" id="path3726-1" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" clip-path="url(#clipPath6265-3-4-4-5)"/>
      <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3728-0" style="display:inline;opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:type="arc" clip-path="url(#clipPath6259-8-81-2-8)"/>
    </ns0:g>
    <ns0:g style="display:inline" id="g4692-3" ns1:label="system-shutdown" transform="matrix(1.333369,0,0,1.333369,604.00453,-317.9473)">
      <ns0:rect width="16" height="16" rx="0.14408804" ry="0.15129246" x="40" y="688" id="rect10837-3-0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none;enable-background:new"/>
      <ns0:path ns2:type="arc" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" id="path3869-2" ns2:cx="48" ns2:cy="696" ns2:rx="7" ns2:ry="7" d="m 51.52343,689.95141 a 7,7 0 0 1 3.233191,7.87837 7,7 0 0 1 -6.766907,5.17021 7,7 0 0 1 -6.751683,-5.19008 7,7 0 0 1 3.25633,-7.86883" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" ns2:start="5.239857" ns2:end="4.1878597" ns2:open="true"/>
      <ns0:path ns1:connector-curvature="0" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="m 48,689 v 5" id="path4710" ns2:nodetypes="cc"/>
    </ns0:g>
    <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:4.00010681;marker:none;enable-background:accumulate" d="m 697.48335,610.6326 -5.00012,5.00014 -5.00015,-5.00014 z" id="rect12003" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
    <ns0:g transform="matrix(0.72370712,0,0,0.72370712,-970.694,430.94511)" id="g17780">
      <ns0:g clip-path="url(#clipPath14882)" ns1:export-ydpi="90" ns1:export-xdpi="90" ns1:export-filename="/home/jimmac/gfx/redhat/redhat-ux/Products/RHEL/RHEL7/video-jingles/tex/overview.png" id="g17782" style="display:inline" transform="matrix(1.6234335,0,0,1.6234335,645.35105,529.77601)">
        <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 239.06066,57.414214 800.87864,0 0,51.485276 c 0,0 -4.0279,-10.606597 -11.0989,-10.96015 L 249,99 c -4.59619,-0.353553 -9.93934,5.5 -9.93934,5.5 z" id="path17784" ns1:connector-curvature="0" ns2:nodetypes="ccccccc"/>
        <ns0:g id="g17786" transform="translate(11,0)">
          <ns0:rect y="58.307991" x="229" height="600" width="800" id="rect17788" style="color:#000000;fill:none;stroke:url(#linearGradient17826);stroke-width:1.38776851;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
          <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" d="m 1028.815,108.766 c 0,-5.89806 -4.7813,-10.6794 -10.6794,-10.6794 l -777.99933,0 c -5.89809,0 -10.6794,4.78134 -10.6794,10.6794" style="fill:none;stroke:#000000;stroke-width:1.09781706px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" id="path17790"/>
        </ns0:g>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g17794" transform="matrix(1.333369,0,0,1.333369,600.00453,608.0695)" ns1:label="audio-volume-medium" style="display:inline">
      <ns0:path ns2:nodetypes="ccccccccc" id="path17796" d="m 20,222 h 2.484375 L 25.453129,219 26,219.0156 v 11 l -0.475297,8.3e-4 L 22.484375,227 H 20 Z" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none" ns1:connector-curvature="0"/>
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" id="rect17798" width="16" height="16" x="20" y="217" ns1:label="audio-volume-high"/>
      <ns0:path clip-path="url(#clipPath6279-7-9-7)" ns2:type="arc" style="display:inline;fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" id="path17800" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" ns2:open="true" ns2:start="5.4977871" ns2:end="0.78539819"/>
      <ns0:path clip-path="url(#clipPath6265-3-4-4-5)" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path17802" style="display:inline;fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:type="arc" ns2:open="true" ns2:start="5.4977871" ns2:end="0.78539819"/>
      <ns0:path clip-path="url(#clipPath6259-8-81-2-8)" ns2:type="arc" style="display:inline;opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" id="path17804" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" ns2:open="true" ns2:start="5.4977871" ns2:end="0.78539819"/>
    </ns0:g>
    <ns0:g transform="matrix(1.333369,0,0,1.333369,600.00453,-19.947301)" ns1:label="system-shutdown" id="g17806" style="display:inline">
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none;enable-background:new" id="rect17808" y="688" x="40" ry="0.15129246" rx="0.14408804" height="16" width="16"/>
      <ns0:path ns2:open="true" ns2:end="4.1878597" ns2:start="5.239857" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" d="m 51.52343,689.95141 a 7,7 0 0 1 3.233191,7.87837 7,7 0 0 1 -6.766907,5.17021 7,7 0 0 1 -6.751683,-5.19008 7,7 0 0 1 3.25633,-7.86883" ns2:ry="7" ns2:rx="7" ns2:cy="696" ns2:cx="48" id="path17810" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" ns2:type="arc"/>
      <ns0:path ns2:nodetypes="cc" id="path17812" d="m 48,689 v 5" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="path17824" d="m 693.48335,908.6326 -5.00012,5.00014 -5.00015,-5.00014 z" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:4.00010681;marker:none;enable-background:accumulate"/>
    <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.39755595;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 381.07806,787.85969 5.62229,5.62229 -5.62229,5.6223 z" id="rect18441" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
    <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="path18444" d="m 463.07806,787.85969 5.62229,5.62229 -5.62229,5.6223 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.39755595;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    <ns0:g transform="matrix(1.3749999,0,0,1.3749999,266.20778,355.98747)" style="display:inline;stroke-width:0.72727281;enable-background:new" ns1:label="network-wired-offline" id="g8415-0">
      <ns0:path ns1:connector-curvature="0" style="color:#bebebe;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:0.35;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#0b0d0d;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" d="m -175,351 v 5 h 2 v 2 h -4.96875 v 3 H -180 v 4.9375 h 5 V 361 h -1.96875 v -2 H -168 v 0.98353 h 1 V 358 h -5 v -2 h 2 v -5 z" transform="translate(421.0002,-173)" id="rect8421-6" ns2:nodetypes="ccccccccccccccccccccc"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="ccccccccccccccccc" id="path3761-2-3-5-4-8-9-8-0-1-7-8-7" d="m 252.0002,188 h 1.375 l 1.125,1.09375 L 255.59395,188 h 1.40625 v 1.46875 l -1.09375,1.0625 1.09375,1.0625 V 193 h -1.4375 l -1.0625,-1.0625 -1.0625,1.0625 h -1.4375 v -1.40625 l 1.0625,-1.0625 -1.0625,-1.0625 z" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#0b0d0d;fill-opacity:1;stroke:none;stroke-width:1.45454562;marker:none"/>
    </ns0:g>
    <ns0:g transform="matrix(1.9999998,0,0,1.9999998,-154.00075,424.00004)" style="display:inline;stroke-width:0.50000006;enable-background:new" ns1:label="network-wired-offline" id="g8415-0-3">
      <ns0:rect y="177" x="241.0002" height="16" width="16" id="rect8417-3" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.50000006;marker:none"/>
      <ns0:path ns1:connector-curvature="0" style="color:#bebebe;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:0.35;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" d="m -175,351 v 5 h 2 v 2 h -4.96875 v 3 H -180 v 4.9375 h 5 V 361 h -1.96875 v -2 H -168 v 0.98353 h 1 V 358 h -5 v -2 h 2 v -5 z" transform="translate(421.0002,-173)" id="rect8421-6-1" ns2:nodetypes="ccccccccccccccccccccc"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="ccccccccccccccccc" id="path3761-2-3-5-4-8-9-8-0-1-7-8-7-5" d="m 252.0002,188 h 1.375 l 1.125,1.09375 L 255.59395,188 h 1.40625 v 1.46875 l -1.09375,1.0625 1.09375,1.0625 V 193 h -1.4375 l -1.0625,-1.0625 -1.0625,1.0625 h -1.4375 v -1.40625 l 1.0625,-1.0625 -1.0625,-1.0625 z" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1.00000012;marker:none"/>
    </ns0:g>
    <ns0:g id="g12704" ns1:label="network-wired-acquiring" style="display:inline;stroke-width:0.5;enable-background:new" transform="matrix(2,0,0,2,-72.000397,423.9437)">
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.5;marker:none" id="rect12706" width="16" height="16" x="241.0002" y="177"/>
      <ns0:rect style="color:#bebebe;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:0.35;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" id="rect12733" width="5.0160389" height="4.9718447" x="240.97597" y="187.98824"/>
      <ns0:rect y="178.02815" x="246.0002" height="4.9718447" width="5.0160389" id="rect12735" style="color:#bebebe;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:0.35;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate"/>
      <ns0:rect style="color:#bebebe;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:0.35;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" id="rect12737" width="5.0160389" height="4.9718447" x="252.0002" y="188.02815"/>
      <ns0:rect style="color:#000000;clip-rule:nonzero;display:block;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#0c0e0e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:new" id="rect11487" width="2.9922597" height="2.9971614" x="243.02184" y="184.04089" rx="0.74806494" ry="0.74806494"/>
      <ns0:rect ry="0.74806494" rx="0.74806494" y="184.04089" x="247.02185" height="2.9971614" width="2.9922597" id="rect11504" style="color:#000000;clip-rule:nonzero;display:block;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#2e3436;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:new"/>
      <ns0:rect style="color:#000000;clip-rule:nonzero;display:block;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#0c0e0e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:new" id="rect11506" width="2.9922597" height="2.9971614" x="247.02185" y="184.04089" rx="0.74806494" ry="0.74806494"/>
      <ns0:rect ry="0.74806494" rx="0.74806494" y="184.04089" x="251.02185" height="2.9971614" width="2.9922597" id="rect11528" style="color:#000000;clip-rule:nonzero;display:block;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#0c0e0e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:new"/>
    </ns0:g>
    <ns0:g style="display:inline;enable-background:new" ns1:label="network-wired" id="g8415" transform="matrix(1.9999997,0,0,1.9999997,2.9996746,424.00005)">
      <ns0:rect y="177" x="241.0002" height="16" width="16" id="rect8417" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none"/>
      <ns0:rect ry="0" y="188" x="241.0002" height="4.9375" width="5.0000014" id="rect8421" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#1a1d1e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate"/>
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#1a1d1e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate" id="rect8425" width="5.0000014" height="5.0000024" x="251.0002" y="188" ry="0"/>
      <ns0:path style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" d="M 2.53125,-8.4687501 V -11.5 H 12.5 v 3.0312499" id="path8427" ns1:connector-curvature="0" transform="translate(241.0002,197)" ns2:nodetypes="cccc"/>
      <ns0:path style="fill:none;stroke:#171a1b;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" d="M 7.5,-11.5 V -15" id="path9198" ns1:connector-curvature="0" transform="translate(241.0002,197)"/>
      <ns0:rect ry="0" y="178" x="246.0002" height="5.0000024" width="5.0000014" id="rect9200" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#1a1d1e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate"/>
    </ns0:g>
    <ns0:g style="display:inline;enable-background:new" ns1:label="network-wired" id="g8415-1" transform="matrix(1.3749998,0,0,1.3749998,263.13713,652.86812)">
      <ns0:rect y="177" x="241.0002" height="16" width="16" id="rect8417-8" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none"/>
      <ns0:rect ry="0" y="188" x="241.0002" height="4.9375" width="5.0000014" id="rect8421-4" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#1a1d1e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate"/>
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#1a1d1e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate" id="rect8425-1" width="5.0000014" height="5.0000024" x="251.0002" y="188" ry="0"/>
      <ns0:path style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" d="M 2.53125,-8.4687501 V -11.5 H 12.5 v 3.0312499" id="path8427-3" ns1:connector-curvature="0" transform="translate(241.0002,197)" ns2:nodetypes="cccc"/>
      <ns0:path style="fill:none;stroke:#171a1b;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" d="M 7.5,-11.5 V -15" id="path9198-9" ns1:connector-curvature="0" transform="translate(241.0002,197)"/>
      <ns0:rect ry="0" y="178" x="246.0002" height="5.0000024" width="5.0000014" id="rect9200-5" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#1a1d1e;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate"/>
    </ns0:g>
  </ns0:g>
</ns0:svg>
