<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="500" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-goa5.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17453" ns4:href="#linearGradient5716" ns1:collect="always"/>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17455" ns4:href="#linearGradient5716" ns1:collect="always"/>
    <ns0:filter color-interpolation-filters="sRGB" ns1:collect="always" x="-0.10291173" width="1.2058235" y="-0.065432459" height="1.1308649" id="filter5601">
      <ns0:feGaussianBlur ns1:collect="always" stdDeviation="0.610872" id="feGaussianBlur5603"/>
    </ns0:filter>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17453-7" ns4:href="#linearGradient5716-4" ns1:collect="always"/>
    <ns0:linearGradient id="linearGradient5716-4">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-1"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-6"/>
    </ns0:linearGradient>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17455-1" ns4:href="#linearGradient5716-4" ns1:collect="always"/>
    <ns0:linearGradient id="linearGradient16929">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop16931"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop16933"/>
    </ns0:linearGradient>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="383.02942" ns1:cy="302.54948" ns1:document-units="px" ns1:current-layer="layer2" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="1484" ns1:window-height="1249" ns1:window-x="355" ns1:window-y="132" ns1:window-maximized="0" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="656" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-540)">
    <ns0:g id="g11020" transform="translate(-35,-141.36217)">
      <ns0:circle transform="translate(2,453.36217)" id="path11014" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;enable-background:accumulate" cx="120" cy="278" r="17"/>
      <ns0:text id="text11016" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan11018" ns2:role="line" style="font-size:14px;line-height:1.25">6</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g style="display:inline" id="g4890" transform="matrix(2.6833333,0,0,2.6833333,-1275.5101,-1072.8539)">
      <ns0:g style="display:inline" id="default-pointer-c" ns1:label="#g5607" transform="matrix(1.0281734,0,0,1.0281734,813.41674,729.17439)">
        <ns0:path ns1:connector-curvature="0" style="opacity:0.6;color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;filter:url(#filter5601);enable-background:accumulate" d="m 27.135224,2.8483222 0,16.4402338 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 27.135224,2.8483222 z" id="path5567" ns2:nodetypes="cccccccc"/>
        <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccccccc" id="path5565" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" style="color:#000000;fill:url(#linearGradient17453-7);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate"/>
        <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:url(#linearGradient17455-1);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path6242" ns2:nodetypes="cccccccc"/>
      </ns0:g>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect4889" width="167.70187" height="168.81989" x="556.96027" y="608.88965"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.47858" y="635.46222" id="text26176"><ns0:tspan ns2:role="line" id="tspan26178" x="610.47858" y="635.46222" style="font-size:5.21739101px;line-height:1.25">Google</ns0:tspan></ns0:text>
      <ns0:text id="text26182" y="642.17023" x="610.47858" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="642.17023" x="610.47858" id="tspan26184" ns2:role="line" style="font-size:4.47205019px;line-height:1.25">maria.johansson@gmail.com</ns0:tspan></ns0:text>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="611.59662" y="666.76648" id="text26186"><ns0:tspan ns2:role="line" id="tspan26188" x="611.59662" y="666.76648" style="font-size:5.21739101px;line-height:1.25">Använd för</ns0:tspan></ns0:text>
      <ns0:text id="text26190" y="666.76648" x="622.40393" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="666.76648" x="622.40393" id="tspan26192" ns2:role="line" style="font-size:5.21739101px;line-height:1.25">E-post</ns0:tspan></ns0:text>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="679.43726" id="text28655"><ns0:tspan ns2:role="line" id="tspan28657" x="622.40393" y="679.43726" style="font-size:5.21739101px;line-height:1.25">Kalender</ns0:tspan></ns0:text>
      <ns0:text id="text28673" y="692.10803" x="622.40393" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="692.10803" x="622.40393" id="tspan28675" ns2:role="line" style="font-size:5.21739101px;line-height:1.25">Kontakter</ns0:tspan></ns0:text>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="704.77881" id="text28691"><ns0:tspan ns2:role="line" id="tspan28693" x="622.40393" y="704.77881" style="font-size:5.21739101px;line-height:1.25">Foto</ns0:tspan></ns0:text>
      <ns0:text id="text28709" y="717.44958" x="622.40393" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="717.44958" x="622.40393" id="tspan28711" ns2:role="line" style="font-size:5.21739101px;line-height:1.25">Filer</ns0:tspan></ns0:text>
      <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect3923-9" width="19.803892" height="10.92049" x="670.62494" y="660.20514" rx="5.4602423" ry="5.4602423"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="path915" cx="684.57684" cy="665.66193" r="4.4139271"/>
      <ns0:path style="opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="path4883" ns2:type="arc" ns2:cx="595.53174" ns2:cy="636.65363" ns2:rx="5.3133016" ns2:ry="5.3133016" ns2:start="0" ns2:end="5.2359878" ns2:open="true" d="m 600.84504,636.65363 a 5.3133016,5.3133016 0 0 1 -3.93812,5.13225 5.3133016,5.3133016 0 0 1 -5.97664,-2.4756 5.3133016,5.3133016 0 0 1 0.84439,-6.41373 5.3133016,5.3133016 0 0 1 6.41372,-0.84438"/>
      <ns0:path style="color:#000000;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:sans-serif;font-variant-ligatures:normal;font-variant-position:normal;font-variant-caps:normal;font-variant-numeric:normal;font-variant-alternates:normal;font-feature-settings:normal;text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;text-decoration-style:solid;text-decoration-color:#000000;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-orientation:mixed;dominant-baseline:auto;baseline-shift:baseline;text-anchor:start;white-space:normal;shape-padding:0;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" d="m 595.9382,635.63421 v 2.53516 h 5.48321 l 0.69267,-1.30041 0.0155,-1.23475 z" id="path4885" ns1:connector-curvature="0" ns2:nodetypes="cccccc"/>
      <ns0:rect ry="5.4602423" rx="5.4602423" y="672.8761" x="670.62494" height="10.92049" width="19.803892" id="rect4891" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
      <ns0:circle r="4.4139271" cy="678.33289" cx="684.57684" id="circle4893" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect ry="5.4602423" rx="5.4602423" y="685.54669" x="670.62494" height="10.92049" width="19.803892" id="rect4899" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
      <ns0:circle r="4.4139271" cy="691.00348" cx="684.57684" id="circle4901" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect4903" width="19.803892" height="10.92049" x="670.62494" y="698.21765" rx="5.4602423" ry="5.4602423"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle4905" cx="684.57684" cy="703.67444" r="4.4139271"/>
      <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect4907" width="19.803892" height="10.92049" x="670.62494" y="710.88824" rx="5.4602423" ry="5.4602423"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle4909" cx="684.57684" cy="716.34503" r="4.4139271"/>
      <ns0:rect ry="5.4602423" rx="5.4602423" y="723.5592" x="670.62494" height="10.92049" width="19.803892" id="rect4911" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
      <ns0:circle r="4.4139271" cy="729.01599" cx="684.57684" id="circle4913" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="730.86591" id="text4917"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" ns2:role="line" id="tspan4915" x="622.40393" y="730.86591">Skriv­ar­e</ns0:tspan></ns0:text>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#c01c28;fill-opacity:1;stroke:none;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect4919" width="54.782524" height="16.397507" x="659.81744" y="750.8772" rx="2.9813664" ry="2.9813664"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.46583843px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.3726708" x="666.71997" y="760.92218" id="text4923"><ns0:tspan ns2:role="line" id="tspan4921" x="666.71997" y="760.92218" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.46583843px;font-family:Cantarell;-inkscape-font-specification:Cantarell;fill:#ffffff;stroke-width:0.3726708">Ta bort konto</ns0:tspan></ns0:text>
    </ns0:g>
  </ns0:g>
</ns0:svg>
