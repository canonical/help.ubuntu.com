<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" height="1000" id="svg10075" version="1.1" width="840" ns2:docname="gs-goa4.svg" ns1:version="0.48.4 r9939">
  <ns0:defs id="defs10077">
    <ns0:linearGradient id="RHEL7" ns3:paint="gradient">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop id="stop11074" offset="0" style="stop-color:#eeedec;stop-opacity:1;"/>
      <ns0:stop id="stop11076" offset="1" style="stop-color:#eeedec;stop-opacity:1"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop id="stop7012" offset="0" style="stop-color:#eeedec;stop-opacity:0;"/>
      <ns0:stop id="stop7014" offset="1" style="stop-color:#eeedec;stop-opacity:0"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(1.1834379,0,0,1.4157524,5.7016703,-219.13426)" gradientUnits="userSpaceOnUse" id="linearGradient7064" x1="-18.33782" x2="713.42853" y1="490.54935" y2="490.54935" ns1:collect="always" ns4:href="#GNOME"/>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient5885" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop id="stop5718" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17441" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop id="stop17445" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop17447" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath24278">
      <ns0:path d="m 0,0 0,2482 2306,0 L 2306,0 0,0 z" id="path24280" ns1:connector-curvature="0"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns2:namedview bordercolor="#666666" borderlayer="true" borderopacity="1.0" fit-margin-bottom="0" fit-margin-left="0" fit-margin-right="0" fit-margin-top="0" height="0px" id="base" pagecolor="#eeeeec" showgrid="false" width="0px" ns1:current-layer="layer3" ns1:cx="-54.723657" ns1:cy="279.56617" ns1:document-units="px" ns1:pageopacity="1" ns1:pageshadow="2" ns1:showpageshadow="false" ns1:snap-bbox="true" ns1:snap-nodes="false" ns1:window-height="1249" ns1:window-maximized="0" ns1:window-width="1484" ns1:window-x="939" ns1:window-y="119" ns1:zoom="0.35355339">
    <ns1:grid empspacing="5" enabled="true" id="grid17504" snapvisiblegridlinesonly="true" type="xygrid" visible="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g id="layer1" transform="translate(0,-492.3622)" ns2:insensitive="true" ns1:groupmode="layer" ns1:label="bg">
    <ns0:rect height="1036" id="background" style="fill:url(#BLANK);" width="866" x="-16" y="475.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g id="layer2" transform="translate(0,-40)" ns1:groupmode="layer" ns1:label="fg">
    <ns0:g id="g11020" transform="translate(-35,-619.36217)">
      <ns0:path d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(2,453.36217)" ns2:cx="120" ns2:cy="278" ns2:rx="17" ns2:ry="17" ns2:type="arc"/>
      <ns0:text id="text11016" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="122.29289" y="736.36218" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan11018" x="122.29289" y="736.36218" ns2:role="line">4</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g id="g24937" transform="translate(17.5,0)">
      <ns0:rect height="411.99997" id="rect17558" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:5.36666679;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="523" x="141" y="105"/>
      <ns0:text id="text12012-1" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="409.45731" y="130.83698" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan12014-2" x="409.45731" y="130.83698" ns2:role="line">Google-konto</ns0:tspan></ns0:text>
      <ns0:rect height="313.93021" id="rect12010-4" rx="0.38461545" ry="0.36744055" style="color:#000000;fill:#eeeeec;stroke:#000000;stroke-width:1.96981525;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="505.19278" x="150.00003" y="150"/>
      <ns0:g id="g17909" transform="translate(73,-471)">
        <ns0:rect height="30.684212" id="rect17494-2" rx="6.1369629" ry="6.1369629" style="color:#000000;fill:none;stroke:#000000;stroke-width:1.99999988;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="96" x="486" y="944"/>
        <ns0:text id="text17496-8" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell" x="533.99988" y="964.00006" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan17498-4" x="533.99988" y="964.00006" ns2:role="line">Avbryt</ns0:tspan></ns0:text>
      </ns0:g>
      <ns0:g clip-path="url(#clipPath24278)" id="g24276" style="fill:#babdb6" transform="matrix(0.125,0,0,-0.125,110.65256,325.93813)">
        <ns0:path d="m 1053.22,1147.46 c 6.96,6.88 7.55,16.45 7.55,21.85 0,21.6 -12.89,55.06 -38.1,55.06 -7.86,0 -16.35,-3.84 -21.15,-9.83 -5.153,-6.34 -6.7,-14.43 -6.7,-22.15 0,-20.05 11.82,-53.34 37.92,-53.34 7.47,0 15.68,3.61 20.48,8.41 z m -8.72,-56.93 -6.94,0.32 c -2.78,0 -19.08,-0.64 -31.78,-4.83 -6.721,-2.39 -26.022,-9.49 -26.022,-30.8 0,-21.31 20.872,-36.49 53.262,-36.49 29,0 44.55,13.8 44.55,32.28 0,15.31 -10.09,23.39 -33.07,39.52 z m 21.42,132.98 c 6.98,-5.68 21.53,-17.63 21.53,-40.42 0,-22.15 -12.63,-32.59 -25.43,-42.54 -3.95,-3.88 -8.5,-8.08 -8.5,-14.67 0,-6.61 4.55,-10.14 7.91,-12.88 l 10.87,-8.39 c 13.32,-11.07 25.46,-21.28 25.46,-41.95 0,-28.05 -27.56,-56.54 -79.6,-56.54 -43.918,0 -65.09,20.64 -65.09,42.89 0,10.72 5.465,25.96 23.321,36.46 18.765,11.37 44.229,12.87 57.799,13.76 -4.18,5.38 -9.06,11.09 -9.06,20.39 0,5.09 1.49,8.08 3.05,11.68 l -9.7,-0.59 c -32.109,0 -50.277,23.63 -50.277,46.98 0,13.75 6.402,29.07 19.402,40.14 17.275,14.09 37.795,16.48 54.165,16.48 l 62.34,0 -19.36,-10.8 -18.83,0" id="path24284" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 913.219,1119.56 c 7.172,9.59 9.078,21.51 9.078,33.16 0,26.39 -12.707,76.55 -50.184,76.55 -9.98,0 -19.972,-3.85 -27.175,-10.16 -11.813,-10.48 -13.879,-23.6 -13.879,-36.46 0,-29.58 14.769,-78.28 51.347,-78.28 11.742,0 23.895,5.68 30.813,15.19 z m -37.793,-24.16 c -48.047,0 -73.75,37.05 -73.75,70.54 0,39.13 32.41,72.62 78.324,72.62 44.375,0 72.113,-34.35 72.113,-70.6 0,-35.28 -27.445,-72.56 -76.687,-72.56" id="path24286" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 749.449,1119.56 c 7.262,9.59 9.012,21.51 9.012,33.16 0,26.39 -12.703,76.55 -50.078,76.55 -9.91,0 -19.992,-3.85 -27.305,-10.16 -11.719,-10.48 -13.836,-23.6 -13.836,-36.46 0,-29.58 14.832,-78.28 51.434,-78.28 11.808,0 23.765,5.68 30.773,15.19 z m -37.824,-24.16 c -48.012,0 -73.777,37.05 -73.777,70.54 0,39.13 32.449,72.62 78.367,72.62 44.39,0 72.14,-34.35 72.14,-70.6 0,-35.28 -27.433,-72.56 -76.73,-72.56" id="path24288" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 614.809,1100.12 -43.379,-10.01 c -17.637,-2.68 -33.496,-5.07 -50.168,-5.07 -83.856,0 -115.703,60.98 -115.703,108.77 0,58.36 45.226,112.4 122.722,112.4 16.391,0 32.184,-2.4 46.442,-6.31 22.793,-6.32 33.445,-14.06 40.086,-18.65 l -25.164,-23.75 -10.657,-2.37 7.578,12.01 c -10.316,9.89 -29.093,28.26 -65.027,28.26 -47.984,0 -84.133,-36.06 -84.133,-88.64 0,-56.49 41.305,-109.72 107.574,-109.72 19.454,0 29.438,3.87 38.571,7.54 l 0,48.36 -45.863,-2.43 24.253,12.99 64.442,0 -7.887,-7.52 -3.058,-4.83 -0.629,-14.44 0,-36.59" id="path24290" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1162.05,1108.67 c -10.08,0.93 -12.14,2.7 -12.14,14.45 l 0,170.11 0.11,1.92 c 1.2,10.56 4.3,12.35 13.71,17.74 l -43.51,0 -22.77,-10.76 23.19,0 0,-0.17 0,0.07 0,-185.54 c 0,-6 -1.15,-6.89 -8.14,-15.92 l 53.77,0 11.19,6.61 c -5.13,0.64 -10.3,0.89 -15.41,1.49" id="path24292" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1257.26,1194.89 c 5.69,2.09 8.73,3.9 8.73,8.05 0,11.89 -13.52,25.72 -29.82,25.72 -12.15,0 -34.77,-9.31 -34.77,-41.52 0,-5.08 0.59,-10.44 0.92,-15.88 l 54.94,23.63 z m 28.33,-88.93 -9.92,-5.4 c -9.97,-4.46 -20.26,-5.68 -29.29,-5.68 -9.65,0 -24.71,0.64 -40.14,11.67 -21.36,14.88 -30.7,40.57 -30.7,62.95 0,46.31 37.99,68.96 69.06,68.96 10.81,0 22.04,-2.71 31.07,-8.34 15.07,-9.86 18.98,-22.73 21.08,-29.57 l -70.81,-28.34 -23.4,-1.81 c 7.62,-37.93 33.63,-59.96 62.22,-59.96 15.39,0 26.58,5.33 36.88,10.39 l -16.05,-14.87" id="path24294" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1314.75,1236.37 0,-19.64 -2.49,0 0,19.64 -6.54,0 0,2.09 15.59,0 0,-2.09 -6.56,0" id="path24296" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1341.89,1216.73 0,19.87 -0.17,0 -6.08,-19.87 -1.94,0 -6.09,19.87 -0.15,0 0,-19.87 -2.2,0 0,21.73 3.76,0 5.65,-17.59 0,0 5.57,17.59 3.76,0 0,-21.73 -2.11,0" id="path24298" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:rect height="34" id="rect24895" style="color:#000000;fill:#cc0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="106" x="538" y="162"/>
      <ns0:text id="text24897" style="font-size:12px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="594" y="183" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24899" x="594" y="183" ns2:role="line">REGISTRERA DIG</ns0:tspan></ns0:text>
      <ns0:text id="text24901" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;font-family:Sans;-inkscape-font-specification:Sans" x="163" y="226" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24903" x="163" y="226" ns2:role="line">Logga in</ns0:tspan></ns0:text>
      <ns0:text id="text24905" style="font-size:13px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;font-family:Sans;-inkscape-font-specification:Sans Bold" x="163" y="259" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24907" x="163" y="259" ns2:role="line">E-post</ns0:tspan></ns0:text>
      <ns0:rect height="35" id="rect24909" rx="0.38461545" ry="0.36744055" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#babdb6;stroke-width:1;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="480" x="164.5" y="265.5"/>
      <ns0:text id="text24911" style="font-size:13px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;font-family:Sans;-inkscape-font-specification:Sans Bold" x="163" y="329" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24913" x="163" y="329" ns2:role="line">Lösenord</ns0:tspan></ns0:text>
      <ns0:rect height="35" id="rect24915" rx="0.38461545" ry="0.36744055" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#babdb6;stroke-width:1;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="480" x="164.5" y="335.5"/>
      <ns0:rect height="34" id="rect24917" style="color:#000000;fill:#729fcf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="106" x="164" y="385"/>
      <ns0:text id="text24919" style="font-size:12px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="218" y="406" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24921" x="218" y="406" ns2:role="line">Logga in</ns0:tspan></ns0:text>
      <ns0:text id="text24923" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;font-family:Sans;-inkscape-font-specification:Sans" x="173" y="287" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24925" x="173" y="287" ns2:role="line">maria.johansson@gmail.com</ns0:tspan></ns0:text>
      <ns0:path d="m 188,294.5 c 0,3.58985 -2.91015,6.5 -6.5,6.5 -3.58985,0 -6.5,-2.91015 -6.5,-6.5 0,-3.58985 2.91015,-6.5 6.5,-6.5 3.58985,0 6.5,2.91015 6.5,6.5 z" id="path24927" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(-1,58)" ns2:cx="181.5" ns2:cy="294.5" ns2:rx="6.5" ns2:ry="6.5" ns2:type="arc"/>
      <ns0:path d="m 188,294.5 c 0,3.58985 -2.91015,6.5 -6.5,6.5 -3.58985,0 -6.5,-2.91015 -6.5,-6.5 0,-3.58985 2.91015,-6.5 6.5,-6.5 3.58985,0 6.5,2.91015 6.5,6.5 z" id="path24929" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(15,58)" ns2:cx="181.5" ns2:cy="294.5" ns2:rx="6.5" ns2:ry="6.5" ns2:type="arc"/>
      <ns0:path d="m 188,294.5 c 0,3.58985 -2.91015,6.5 -6.5,6.5 -3.58985,0 -6.5,-2.91015 -6.5,-6.5 0,-3.58985 2.91015,-6.5 6.5,-6.5 3.58985,0 6.5,2.91015 6.5,6.5 z" id="path24931" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(31,58)" ns2:cx="181.5" ns2:cy="294.5" ns2:rx="6.5" ns2:ry="6.5" ns2:type="arc"/>
      <ns0:path d="m 188,294.5 c 0,3.58985 -2.91015,6.5 -6.5,6.5 -3.58985,0 -6.5,-2.91015 -6.5,-6.5 0,-3.58985 2.91015,-6.5 6.5,-6.5 3.58985,0 6.5,2.91015 6.5,6.5 z" id="path24933" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(47,58)" ns2:cx="181.5" ns2:cy="294.5" ns2:rx="6.5" ns2:ry="6.5" ns2:type="arc"/>
      <ns0:path d="m 188,294.5 c 0,3.58985 -2.91015,6.5 -6.5,6.5 -3.58985,0 -6.5,-2.91015 -6.5,-6.5 0,-3.58985 2.91015,-6.5 6.5,-6.5 3.58985,0 6.5,2.91015 6.5,6.5 z" id="path24935" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(63,58)" ns2:cx="181.5" ns2:cy="294.5" ns2:rx="6.5" ns2:ry="6.5" ns2:type="arc"/>
    </ns0:g>
    <ns0:g id="g24977" transform="translate(17.5,460)">
      <ns0:rect height="411.99997" id="rect24979" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:5.36666679;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="523" x="141" y="105"/>
      <ns0:text id="text24981" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="409.45731" y="130.83698" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24983" x="409.45731" y="130.83698" ns2:role="line">Google-konto</ns0:tspan></ns0:text>
      <ns0:rect height="313.93021" id="rect24985" rx="0.38461545" ry="0.36744055" style="color:#000000;fill:#eeeeec;stroke:#000000;stroke-width:1.96981525;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="505.19278" x="150.00003" y="150"/>
      <ns0:g id="g24987" transform="translate(73,-471)">
        <ns0:rect height="30.684212" id="rect24989" rx="6.1369629" ry="6.1369629" style="color:#000000;fill:none;stroke:#000000;stroke-width:1.99999988;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="96" x="486" y="944"/>
        <ns0:text id="text24991" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell" x="532.99988" y="964.00006" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan24993" x="532.99988" y="964.00006" ns2:role="line">Avbryt</ns0:tspan></ns0:text>
      </ns0:g>
      <ns0:g clip-path="url(#clipPath24278)" id="g24995" style="fill:#babdb6" transform="matrix(0.125,0,0,-0.125,110.65256,325.93813)">
        <ns0:path d="m 1053.22,1147.46 c 6.96,6.88 7.55,16.45 7.55,21.85 0,21.6 -12.89,55.06 -38.1,55.06 -7.86,0 -16.35,-3.84 -21.15,-9.83 -5.153,-6.34 -6.7,-14.43 -6.7,-22.15 0,-20.05 11.82,-53.34 37.92,-53.34 7.47,0 15.68,3.61 20.48,8.41 z m -8.72,-56.93 -6.94,0.32 c -2.78,0 -19.08,-0.64 -31.78,-4.83 -6.721,-2.39 -26.022,-9.49 -26.022,-30.8 0,-21.31 20.872,-36.49 53.262,-36.49 29,0 44.55,13.8 44.55,32.28 0,15.31 -10.09,23.39 -33.07,39.52 z m 21.42,132.98 c 6.98,-5.68 21.53,-17.63 21.53,-40.42 0,-22.15 -12.63,-32.59 -25.43,-42.54 -3.95,-3.88 -8.5,-8.08 -8.5,-14.67 0,-6.61 4.55,-10.14 7.91,-12.88 l 10.87,-8.39 c 13.32,-11.07 25.46,-21.28 25.46,-41.95 0,-28.05 -27.56,-56.54 -79.6,-56.54 -43.918,0 -65.09,20.64 -65.09,42.89 0,10.72 5.465,25.96 23.321,36.46 18.765,11.37 44.229,12.87 57.799,13.76 -4.18,5.38 -9.06,11.09 -9.06,20.39 0,5.09 1.49,8.08 3.05,11.68 l -9.7,-0.59 c -32.109,0 -50.277,23.63 -50.277,46.98 0,13.75 6.402,29.07 19.402,40.14 17.275,14.09 37.795,16.48 54.165,16.48 l 62.34,0 -19.36,-10.8 -18.83,0" id="path24997" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 913.219,1119.56 c 7.172,9.59 9.078,21.51 9.078,33.16 0,26.39 -12.707,76.55 -50.184,76.55 -9.98,0 -19.972,-3.85 -27.175,-10.16 -11.813,-10.48 -13.879,-23.6 -13.879,-36.46 0,-29.58 14.769,-78.28 51.347,-78.28 11.742,0 23.895,5.68 30.813,15.19 z m -37.793,-24.16 c -48.047,0 -73.75,37.05 -73.75,70.54 0,39.13 32.41,72.62 78.324,72.62 44.375,0 72.113,-34.35 72.113,-70.6 0,-35.28 -27.445,-72.56 -76.687,-72.56" id="path24999" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 749.449,1119.56 c 7.262,9.59 9.012,21.51 9.012,33.16 0,26.39 -12.703,76.55 -50.078,76.55 -9.91,0 -19.992,-3.85 -27.305,-10.16 -11.719,-10.48 -13.836,-23.6 -13.836,-36.46 0,-29.58 14.832,-78.28 51.434,-78.28 11.808,0 23.765,5.68 30.773,15.19 z m -37.824,-24.16 c -48.012,0 -73.777,37.05 -73.777,70.54 0,39.13 32.449,72.62 78.367,72.62 44.39,0 72.14,-34.35 72.14,-70.6 0,-35.28 -27.433,-72.56 -76.73,-72.56" id="path25001" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 614.809,1100.12 -43.379,-10.01 c -17.637,-2.68 -33.496,-5.07 -50.168,-5.07 -83.856,0 -115.703,60.98 -115.703,108.77 0,58.36 45.226,112.4 122.722,112.4 16.391,0 32.184,-2.4 46.442,-6.31 22.793,-6.32 33.445,-14.06 40.086,-18.65 l -25.164,-23.75 -10.657,-2.37 7.578,12.01 c -10.316,9.89 -29.093,28.26 -65.027,28.26 -47.984,0 -84.133,-36.06 -84.133,-88.64 0,-56.49 41.305,-109.72 107.574,-109.72 19.454,0 29.438,3.87 38.571,7.54 l 0,48.36 -45.863,-2.43 24.253,12.99 64.442,0 -7.887,-7.52 -3.058,-4.83 -0.629,-14.44 0,-36.59" id="path25003" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1162.05,1108.67 c -10.08,0.93 -12.14,2.7 -12.14,14.45 l 0,170.11 0.11,1.92 c 1.2,10.56 4.3,12.35 13.71,17.74 l -43.51,0 -22.77,-10.76 23.19,0 0,-0.17 0,0.07 0,-185.54 c 0,-6 -1.15,-6.89 -8.14,-15.92 l 53.77,0 11.19,6.61 c -5.13,0.64 -10.3,0.89 -15.41,1.49" id="path25005" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1257.26,1194.89 c 5.69,2.09 8.73,3.9 8.73,8.05 0,11.89 -13.52,25.72 -29.82,25.72 -12.15,0 -34.77,-9.31 -34.77,-41.52 0,-5.08 0.59,-10.44 0.92,-15.88 l 54.94,23.63 z m 28.33,-88.93 -9.92,-5.4 c -9.97,-4.46 -20.26,-5.68 -29.29,-5.68 -9.65,0 -24.71,0.64 -40.14,11.67 -21.36,14.88 -30.7,40.57 -30.7,62.95 0,46.31 37.99,68.96 69.06,68.96 10.81,0 22.04,-2.71 31.07,-8.34 15.07,-9.86 18.98,-22.73 21.08,-29.57 l -70.81,-28.34 -23.4,-1.81 c 7.62,-37.93 33.63,-59.96 62.22,-59.96 15.39,0 26.58,5.33 36.88,10.39 l -16.05,-14.87" id="path25007" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1314.75,1236.37 0,-19.64 -2.49,0 0,19.64 -6.54,0 0,2.09 15.59,0 0,-2.09 -6.56,0" id="path25009" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="m 1341.89,1216.73 0,19.87 -0.17,0 -6.08,-19.87 -1.94,0 -6.09,19.87 -0.15,0 0,-19.87 -2.2,0 0,21.73 3.76,0 5.65,-17.59 0,0 5.57,17.59 3.76,0 0,-21.73 -2.11,0" id="path25011" style="fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:rect height="34" id="rect25035" style="color:#000000;fill:#729fcf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="179" x="164" y="219"/>
      <ns0:text id="text25037" style="font-size:12px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="254" y="240" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan25039" x="254" y="240" ns2:role="line">Bevilja åtkomst</ns0:tspan></ns0:text>
      <ns0:rect height="16" id="rect25076" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="451" x="164" y="273"/>
      <ns0:rect height="16" id="rect25078" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="274" x="164" y="298"/>
      <ns0:g id="g25068" transform="translate(189,-166)">
        <ns0:rect height="34" id="rect25070" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="161" x="164" y="385"/>
        <ns0:text id="text25072" style="font-size:12px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#2e3436;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="247" y="406" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan25074" x="247" y="406" ns2:role="line">Förbjud tillträde</ns0:tspan></ns0:text>
      </ns0:g>
      <ns0:rect height="16" id="rect25085" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="119" x="164" y="337"/>
      <ns0:rect height="16" id="rect25087" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="95" x="164" y="362"/>
      <ns0:rect height="16" id="rect25089" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="119" x="164" y="387"/>
      <ns0:rect height="16" id="rect25091" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="95" x="164" y="412"/>
      <ns0:rect height="311" id="rect25093" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="16" x="638.5" y="151"/>
      <ns0:rect height="203" id="rect25095" rx="4.1756759" ry="4.1756759" style="color:#000000;fill:#888a85;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="8.3513517" x="642.5" y="154"/>
    </ns0:g>
    <ns0:g id="g25055" transform="translate(-35,-159.36217)">
      <ns0:path d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" id="path25057" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(2,453.36217)" ns2:cx="120" ns2:cy="278" ns2:rx="17" ns2:ry="17" ns2:type="arc"/>
      <ns0:text id="text25059" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="122.29289" y="736.36218" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan25061" x="122.29289" y="736.36218" ns2:role="line">5</ns0:tspan></ns0:text>
    </ns0:g>
  </ns0:g>
  <ns0:g id="layer3" style="display:none" ns1:groupmode="layer" ns1:label="stuff">
    <ns0:text id="text17640" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="-218.54269" y="669.83698" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan17642" x="-218.54269" y="669.83698" ns2:role="line">Google</ns0:tspan></ns0:text>
    <ns0:text id="text17893" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="-218.54269" y="709.83698" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan17895" x="-218.54269" y="709.83698" ns2:role="line">Facebook</ns0:tspan></ns0:text>
    <ns0:text id="text17897" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="-218.54269" y="749.83698" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan17899" x="-218.54269" y="749.83698" ns2:role="line">Windows Live</ns0:tspan></ns0:text>
    <ns0:text id="text17901" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="-218.54269" y="789.83698" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan17903" x="-218.54269" y="789.83698" ns2:role="line">Microsoft Exchange</ns0:tspan></ns0:text>
    <ns0:text id="text17905" style="font-size:14px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;display:inline;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" x="-218.54269" y="829.83698" ns2:linespacing="125%" xml:space="preserve"><ns0:tspan id="tspan17907" x="-218.54269" y="829.83698" ns2:role="line">Företagsinloggning (Kerberos)</ns0:tspan></ns0:text>
    <ns0:g id="g3922" style="display:inline" transform="matrix(2,0,0,2,-302,333)" ns1:label="account-facebook">
      <ns0:rect height="16" id="rect2941" style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" transform="matrix(0,-1,1,0,0,0)" width="16" x="-194" y="20" ns1:label="audio-volume-high"/>
      <ns0:path d="M 22.116732,178 C 20.946094,178 20,178.94979 20,180.125 l 0,11.75 c 0,1.17521 0.946094,2.125 2.116732,2.125 l 6.910506,0 0,-6 -0.99611,0 0,-2 0.99611,0 0,-1.0625 c 0,-1.84445 1.374066,-2.88912 3.175096,-2.9375 l 1.77432,0 0,2 -1.089494,0 c -0.625856,0 -0.902724,0.22291 -0.902724,0.90625 l 0,1.09375 1.712062,0 -0.217898,2 -1.494164,0 0,6 1.898832,0 C 35.053906,194 36,193.05021 36,191.875 l 0,-11.75 C 36,178.94979 35.053906,178 33.883268,178 z" id="rect14063" style="color:#000000;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:nodetypes="sssscccccscccsscccccsssss" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:path d="m -252.93756,649.01715 -3.56249,-0.016 c -2.51115,1.30826 -2.88681,4.57261 -2.06249,7.56248 1.08953,3.95154 3.26699,6.72334 6.18748,5.81248 4.0738,-1.27088 4.19302,-4.59783 2.93749,-8.49998 -0.66404,-2.06383 -1.89568,-3.7267 -3.49999,-4.85936 z m 9.93747,6.17186 c 0,1.75946 -0.71594,3.26127 -1.5,4.43749 l 0,0.0624 -0.1874,0.125 c 0,0 -0.50952,0.59837 -1.12499,1.18749 -0.61462,0.58922 -1.5625,1.375 -1.5625,1.375 -0.7713,0.57968 -1.1875,1.34601 -1.1875,2.18749 0,0.84434 0.53654,1.6075 1.3125,2.18749 0,0 1.5736,0.96414 2.43749,1.6875 0.86354,0.7238 1.875,1.68749 1.875,1.68749 1.16965,1.09974 1.93749,2.8523 1.93749,4.81249 0,1.68819 -0.5353,3.21907 -1.43749,4.31249 l -1.375,1.74999 8.56247,0 c 2.34128,0 4.24999,-1.89957 4.24999,-4.24999 l 0,-23.49992 c 0,-2.35042 -1.90871,-4.24999 -4.24999,-4.24999 -1.14773,-0.014 -3.64297,0.004 -3.64297,0.004 l -0.031,1.97129 -5.13194,0.57558 c 0.7509,1.3041 1.03662,2.60573 1.05596,3.63721 z m -19.99994,4.87499 0,11.24996 c 3.47287,-2.32521 9.68747,-2.37499 9.68747,-2.37499 0,0 0.027,-0.0372 0,-0.0624 -2.49155,-1.91534 -1.4375,-4.12509 -1.4375,-4.12509 -3.8524,0.3282 -5.61338,-1.10972 -8.24997,-4.68748 z m 10.12497,11.06246 c -3.46111,0.1948 -7.91464,1.6274 -7.99998,5.06249 0,2.05473 1.33766,3.91718 3.24999,4.74998 0,0 0.0688,0.0442 0.125,0.0624 l 0.0624,0 9.06247,0 c 0,0 0.0212,-0.0894 0.0624,-0.125 4.90245,-4.33881 1.20038,-6.85438 -2.99999,-9.68747 -0.0758,-0.0504 -0.1874,-0.0624 -0.1874,-0.0624 -0.43799,-0.0208 -0.88055,-0.0278 -1.37499,0 z" id="path14750" style="color:#000000;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:nodetypes="ccccscscccccscccsccssscccccsccccsccccccccsccc" ns1:connector-curvature="0"/>
  </ns0:g>
</ns0:svg>
