<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Filer, mappar och sökning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Filer, mappar och sökning</span></h1></div>
<div class="region">
<div class="contents">
<div class="media media-image floatend if-if if__not-target-mobile"><div class="inner"><img src="figures/nautilus.png" class="media media-block" alt="Filhanteraren Nautilus"></div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Vanliga åtgärder</span></h2></div>
<div class="region"><ul>
<li class="links "><a class="bold" href="files-browse.html" title="Bläddra bland filer och mappar">Bläddra bland filer och mappar</a></li>
<li class="links "><a class="bold" href="files-rename.html" title="Byt namn på en fil eller mapp">Byt namn på en fil eller mapp</a></li>
<li class="links "><a class="bold" href="files-preview.html" title="Förhandsgranska filer och mappar">Förhandsgranska filer och mappar</a></li>
<li class="links "><a class="bold" href="files-copy.html" title="Kopiera eller flytta filer och mappar">Kopiera eller flytta filer och mappar</a></li>
<li class="links "><a class="bold" href="files-sort.html" title="Sortera filer och mappar">Sortera filer och mappar</a></li>
<li class="links "><a class="bold" href="files-search.html" title="Sök efter filer">Sök efter filer</a></li>
<li class="links "><a class="bold" href="files-delete.html" title="Ta bort filer och mappar">Ta bort filer och mappar</a></li>
</ul></div>
</div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Fler ämnen</span></h2></div>
<div class="region"><ul>
<li class="links "><a class="bold" href="nautilus-connect.html" title="Bläddra bland filer på en server eller nätverksdelning">Bläddra bland filer på en server eller nätverksdelning</a></li>
<li class="links "><a class="bold" href="files-share.html" title="Dela ut och överför filer">Dela ut och överför filer</a></li>
<li class="links "><a class="bold" href="nautilus-file-properties-basic.html" title="Filegenskaper">Filegenskaper</a></li>
<li class="links "><a class="bold" href="files-lost.html" title="Hitta en borttappad fil">Hitta en borttappad fil</a></li>
<li class="links "><a class="bold" href="files-disc-write.html" title="Skriv filer till en cd- eller dvd-skiva">Skriv filer till en cd- eller dvd-skiva</a></li>
<li class="links "><a class="bold" href="files-recover.html" title="Återställ en fil från Papperskorgen">Återställ en fil från Papperskorgen</a></li>
<li class="links "><a class="bold" href="files-open.html" title="Öppna filer med andra program">Öppna filer med andra program</a></li>
<li class="links "><a class="bold" href="nautilus-prefs.html" title="Inställningar för filhanterare">Inställningar för filhanterare</a></li>
</ul></div>
</div></div>
</div>
<div id="removable" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Flyttbara enheter och externa diskar</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="files-removedrive.html" title="Säker borttagning av extern enhet"><span class="title">Säker borttagning av extern enhet</span><span class="linkdiv-dash"> — </span><span class="desc">Mata ut eller avmontera en USB-enhet, CD-/DVD-skiva, eller en annan enhet.</span></a></div></div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="files-autorun.html" title="Öppna program för enheter eller skivor"><span class="title">Öppna program för enheter eller skivor</span><span class="linkdiv-dash"> — </span><span class="desc">Kör automatiskt program för CD- och DVD-skivor, kameror, musikspelare, och andra enheter och media.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="backup" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Säkerhetskopiering</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="backup-frequency.html" title="Frekvens för säkerhetskopiering"><span class="title">Frekvens för säkerhetskopiering</span><span class="linkdiv-dash"> — </span><span class="desc">Få tips om hur ofta du bör ta säkerhetskopior för att se till att dina filer är säkra.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="backup-check.html" title="Kontrollera din säkerhetskopia"><span class="title">Kontrollera din säkerhetskopia</span><span class="linkdiv-dash"> — </span><span class="desc">Kontrollera att din säkerhetskopiering lyckades.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="backup-why.html" title="Säkerhetskopiera dina viktiga filer"><span class="title">Säkerhetskopiera dina viktiga filer</span><span class="linkdiv-dash"> — </span><span class="desc">Varför, vad, var, och hur man säkerhetskopierar.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="backup-thinkabout.html" title="Var hittar jag filerna jag vill säkerhetskopiera?"><span class="title">Var hittar jag filerna jag vill säkerhetskopiera?</span><span class="linkdiv-dash"> — </span><span class="desc">En lista över mappar där du kan hitta dokument, filer och inställningar som du kan vilja kopiera.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="backup-restore.html" title="Återställ en säkerhetskopia"><span class="title">Återställ en säkerhetskopia</span><span class="linkdiv-dash"> — </span><span class="desc">Få tillbaka dina filer från en säkerhetskopia.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="documents" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Dokument</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="documents.html" title="Dokument"><span class="title">Dokument</span><span class="linkdiv-dash"> — </span><span class="desc">Organisera dokumenten som lagras lokalt på din dator eller som skapats på internet.</span></a></div></div>
<div class="links-twocolumn"></div>
</div></div></div></div></div>
</div></div>
<div id="faq" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Tips och frågor</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="nautilus-file-properties-permissions.html" title="Ange filrättigheter"><span class="title">Ange filrättigheter</span><span class="linkdiv-dash"> — </span><span class="desc">Styr vem som kan visa och redigera dina filer och mappar.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-hidden.html" title="Dölj en fil"><span class="title">Dölj en fil</span><span class="linkdiv-dash"> — </span><span class="desc">Gör en fil osynlig, så att du inte kan se den i filhanteraren.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-templates.html" title="Mallar för vanligt förekommande dokumenttyper"><span class="title">Mallar för vanligt förekommande dokumenttyper</span><span class="linkdiv-dash"> — </span><span class="desc">Skapa snabbt nya dokument från egna filmallar.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="files-select.html" title="Markera filer efter mönster"><span class="title">Markera filer efter mönster</span><span class="linkdiv-dash"> — </span><span class="desc">Tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>S</kbd></span></span> för att välja flera filer med liknande namn.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="nautilus-bookmarks-edit.html" title="Redigera mappbokmärken"><span class="title">Redigera mappbokmärken</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till, ta bort och byt namn på bokmärken i filhanteraren.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-tilde.html" title='Vad är en fil med ett "~" i slutet av filnamnet?'><span class="title">Vad är en fil med ett "~" i slutet av filnamnet?</span><span class="linkdiv-dash"> — </span><span class="desc">Detta är säkerhetskopior. De är dolda som standard.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
