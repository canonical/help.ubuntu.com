<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Byt namn på en fil eller mapp</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Byt namn på en fil eller mapp</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan använda filhanteraren för att byta namn på en fil eller mapp.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">För att byta namn på en fil eller mapp:</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Högerklicka på objektet och välj <span class="gui">Byt namn</span> eller markera filen och tryck på <span class="key"><kbd>F2</kbd></span>.</p></li>
<li class="steps"><p class="p">Ange det nya namnet och tryck på <span class="key"><kbd>Retur</kbd></span>.</p></li>
</ol></div>
</div></div>
<p class="p">Du kan också byta namn på en fil från fönstret<span class="link"><a href="nautilus-file-properties-basic.html" title="Filegenskaper">egenskaper</a></span>.</p>
<p class="p">När du döper om en fil markeras bara den första delen av filnamnet, inte filändelsen (biten efter "."). Filändelsen berättar vanligtvis vilken filtyp det är (<span class="file">fil.pdf</span> t.ex. är ett PDF-dokument), och du vill i regel inte ändra den. Om du ändå behöver ändra filändelsen också, markera hela filnamnet manuellt och ändra det.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du döpte om fel fil, eller gav filen ett felaktigt namn, kan du ångra namnbytet. För att backa åtgärden och återställa det tidigare namnet, klicka omedelbart på <span class="gui">Redigera</span> i menyraden och välj <span class="gui">Ångra namnbyte</span>.</p></div></div></div></div>
</div>
<div id="valid-chars" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Giltiga tecken för filnamn</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan använda vilka tecken som helst förutom <span class="key"><kbd>/</kbd></span> (snedstreck) i filnamn. Vissa enheter använder tyvärr ett <span class="em">filsystem</span> som är mer restriktivt vad gäller filnamn. Därför är det god sed att undvika följande tecken i dina filnamn: <span class="key"><kbd>|</kbd></span>, <span class="key"><kbd>\</kbd></span>, <span class="key"><kbd>?</kbd></span>, <span class="key"><kbd>*</kbd></span>, <span class="key"><kbd>&lt;</kbd></span>, <span class="key"><kbd>"</kbd></span>, <span class="key"><kbd>:</kbd></span>, <span class="key"><kbd>&gt;</kbd></span>, <span class="key"><kbd>/</kbd></span>.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du använder filnamn som har en <span class="key"><kbd>.</kbd></span> som första tecken kommer filen bli <span class="link"><a href="files-hidden.html" title="Dölj en fil">dold</a></span> när du försöker visa den i filhanteraren.</p></div></div></div></div>
</div></div>
</div></div>
<div id="common-probs" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Vanliga problem</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Filnamnet används redan</dt>
<dd class="terms">
<p class="p">Du får inte ha två filer eller mappar med samma namn i samma mapp. Om du försöker döpa om en fil till ett namn som redan finns i mappen du arbetar i kommer filhanteraren inte tillåta det.</p>
<p class="p">Fil- och mappnamn gör skillnad på stor och liten bokstav, så filnamnet <span class="file">Fil.txt</span> är inte samma som <span class="file">FIL.txt</span>. Det är tillåtet att använda sådana variationer av filnamn, men det rekommenderas inte.</p>
</dd>
<dt class="terms">Filnamnet är för långt</dt>
<dd class="terms"><p class="p">I vissa filsystem får inte filnamn bestå av fler än 255 tecken. Gränsen på 255 tecken räknar både filnamnet och sökvägen till filen (t.ex. <span class="file">/home/vanja/Dokument/arbete/business-proposals/...</span>), så du bör undvika långa fil- och mappnamn närhelst du kan.</p></dd>
<dt class="terms">Alternativet att byta namn är inaktiverat</dt>
<dd class="terms"><p class="p">Om <span class="gui">Byt namn</span> är blockerat har du inte tillstånd att döpa om filen. Du bör vara försiktig när du försöker döpa om sådana filer, eftersom systemet kan bli instabilt om vissa skydda filer döps om. Se link xref="nautilus-file-properties-permissions"/&gt; för mer information.</p></dd>
</dl></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer eller kataloger">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
