<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Connect to a wireless network</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Connect to a wireless network</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">If you have a wireless-enabled computer, you can connect to a wireless network that is within range to get access to the internet, view shared files on the network, and so on.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">If you have a wireless hardware switch on your computer, make sure that it is turned on.</p></li>
<li class="steps">
<p class="p">Click the <span class="gui">network menu</span> in the <span class="gui">menu bar</span>, and click the name of the network you want to connect to.</p>
<p class="p">If the name of the network isn't in the list, select <span class="gui">More Networks</span> to see if the network is further down the list. If you still don't see the network, you may be out of range or the network <span class="link"><a href="net-wireless-hidden.html" title="Connect to a hidden wireless network">might be hidden</a></span>.</p>
</li>
<li class="steps">
<p class="p">If the network is protected by a password (<span class="link"><a href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?">encryption key</a></span>), enter the password when prompted and click <span class="gui">Connect</span>.</p>
<p class="p">If you do not know the key, it may be written on the underside of the wireless router or base station, in its instruction manual, or you may have to ask the person who administers the wireless network.</p>
</li>
<li class="steps"><p class="p">The network icon will change appearance as the computer attempts to connect to the network.</p></li>
<li class="steps"><p class="p">If the connection is successful, the icon will change to a dot with several bars above it. More bars indicate a stronger connection to the network. If there aren't many bars, the connection is weak and might not be very reliable.</p></li>
</ol></div></div></div>
<p class="p">If the connection is not successful, you <span class="link"><a href="net-wireless-noconnection.html" title="I've entered the correct password, but I still can't connect">may be asked for your password again</a></span> or it might just tell you that the connection has been disconnected. There are a number of things that could have caused this to happen. You could have entered the wrong password, the wireless signal could be too weak, or your computer's wireless card might have a problem, for example. See <span class="link"><a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a></span> for more help.</p>
<p class="p">A stronger connection to a wireless network does not necessarily mean that you have a faster internet connection, or that you will have faster download speeds. The wireless connection connects your computer to the <span class="em">device which provides the internet connection</span> (like a router or modem), but the two connections are actually different, and so will run at different speeds.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a><span class="desc"> — 
      <span class="link"><a href="net-wireless-connect.html" title="Connect to a wireless network">Connect to wifi</a></span>,
      <span class="link"><a href="net-wireless-hidden.html" title="Connect to a hidden wireless network">Hidden networks</a></span>,
      <span class="link"><a href="net-wireless-edit-connection.html" title="Redigera en trådlös anslutning">Edit connection settings</a></span>,
      <span class="link"><a href="net-wireless-disconnecting.html" title="Why does my wireless network keep disconnecting?">Disconnecting</a></span>…
    </span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="net-wireless-noconnection.html" title="I've entered the correct password, but I still can't connect">I've entered the correct password, but I still can't connect</a><span class="desc"> — Double-check the password, try using the pass key instead of the password, turn the wireless card off and on again…</span>
</li>
<li class="links ">
<a href="net-wireless-disconnecting.html" title="Why does my wireless network keep disconnecting?">Why does my wireless network keep disconnecting?</a><span class="desc"> — You might have low signal, or the network might not be letting you connect properly.</span>
</li>
<li class="links ">
<a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a><span class="desc"> — Identify and fix problems with wireless connections</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
