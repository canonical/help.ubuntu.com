<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="468" id="svg1525" version="1.1" ns1:version="0.48.4 r9939" ns2:docname="gs-thumb-launching-apps.svg" ns1:export-filename="/home/jimmac/src/cvs/gnome/gnome-getting-started-docs/getting-started/C/figures/windows-and-workspaces.png" ns1:export-xdpi="90" ns1:export-ydpi="90">
  <ns2:namedview id="base" pagecolor="#ffffff" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="0.0" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="738.77767" ns1:cy="283.00167" ns1:document-units="px" ns1:current-layer="layer3" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="2560" ns1:window-height="1401" ns1:window-x="2560" ns1:window-y="0" ns1:window-maximized="1">
    <ns1:grid type="xygrid" id="grid6208"/>
  </ns2:namedview>
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns1:collect="always" id="linearGradient8346">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop8348"/>
      <ns0:stop style="stop-color:#ffffff;stop-opacity:1" offset="1" id="stop8350"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient3962-1-1-9-5-4-2-1" id="radialGradient17454" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1.3341939,0,0,1.3304716,91.10644,199.8237)" cx="18.247644" cy="15.716079" fx="18.247644" fy="15.716079" r="29.993349"/>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2-1">
      <ns0:stop id="stop3964-5-0-1-9-6-6-6" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6-3" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4-5" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7-6"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3-0" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient10586-8-2-5-1-6-0" id="linearGradient17456" gradientUnits="userSpaceOnUse" gradientTransform="matrix(0.24989036,0,0,0.250888,92.6666,202.07506)" x1="145.16281" y1="-41.407383" x2="144.42656" y2="46.077827"/>
    <ns0:linearGradient id="linearGradient10586-8-2-5-1-6-0" ns1:collect="always">
      <ns0:stop id="stop10588-8-7-5-8-3-4" offset="0" style="stop-color: rgb(172, 197, 237); stop-opacity: 1;"/>
      <ns0:stop id="stop10590-3-6-5-8-3-9" offset="1" style="stop-color: rgb(25, 59, 110); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17368-69" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:linearGradient id="linearGradient6868-5-7-5-4-3-8" ns1:collect="always">
      <ns0:stop id="stop6870-84-7-0-1-8-4" offset="0" style="stop-color: rgb(0, 0, 0); stop-opacity: 1;"/>
      <ns0:stop id="stop6872-0-5-0-7-1-5" offset="1" style="stop-color: rgb(0, 0, 0); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17366-7" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17364" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17374-8" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17372-7" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17370" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17380-2" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17378-0" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17376" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17386-08" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17384-5" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17382" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17392-3" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17390-6" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17388" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17398-2" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17396-0" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17394" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17404-3" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17402-4" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17400" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17410-8" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17408-3" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17406" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17416-8" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17414-5" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-8" id="radialGradient17412" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient10599-4-0-8-1-6" id="radialGradient17418" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1.96261,0,0,1.09426,-74.6625,-21.1211)" cx="77.5625" cy="152.51079" fx="77.5625" fy="152.51079" r="13.03125"/>
    <ns0:linearGradient id="linearGradient10599-4-0-8-1-6" ns1:collect="always">
      <ns0:stop id="stop10601-9-3-6-7-5-5" offset="0" style="stop-color: rgb(255, 255, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop10603-3-0-1-5-1" offset="1" style="stop-color: rgb(255, 255, 255); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:filter color-interpolation-filters="sRGB" id="filter10631-9-5-7-4-7" ns1:collect="always">
      <ns0:feGaussianBlur id="feGaussianBlur10633-6-0-3-5-7" stdDeviation="0.5906498" ns1:collect="always"/>
    </ns0:filter>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient3962-1-1-9-5-4-2-0" id="radialGradient17454-5" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1.3341939,0,0,1.3304716,251.10644,532.18588)" cx="18.247644" cy="15.716079" fx="18.247644" fy="15.716079" r="29.993349"/>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2-0">
      <ns0:stop id="stop3964-5-0-1-9-6-6-34" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6-4" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7-0"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3-6" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient10586-8-2-5-1-6-0-1" id="linearGradient17456-9" gradientUnits="userSpaceOnUse" gradientTransform="matrix(0.24989036,0,0,0.250888,252.6666,534.43724)" x1="145.16281" y1="-41.407383" x2="144.42656" y2="46.077827"/>
    <ns0:linearGradient id="linearGradient10586-8-2-5-1-6-0-1" ns1:collect="always">
      <ns0:stop id="stop10588-8-7-5-8-3-4-7" offset="0" style="stop-color: rgb(172, 197, 237); stop-opacity: 1;"/>
      <ns0:stop id="stop10590-3-6-5-8-3-9-2" offset="1" style="stop-color: rgb(25, 59, 110); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30900" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:linearGradient id="linearGradient6868-5-7-5-4-3-2" ns1:collect="always">
      <ns0:stop id="stop6870-84-7-0-1-8-0" offset="0" style="stop-color: rgb(0, 0, 0); stop-opacity: 1;"/>
      <ns0:stop id="stop6872-0-5-0-7-1-9" offset="1" style="stop-color: rgb(0, 0, 0); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30898" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17364-2" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30904" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30902" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17370-0" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30908" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30906" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17376-6" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30912" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30910" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17382-0" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30916" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30914" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17388-62" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30920" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30918" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17394-9" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30924" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30922" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17400-9" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30928" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30926" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17406-0" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30932" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient30930" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3-2" id="radialGradient17412-86" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient10599-4-0-8-1-6-9" id="radialGradient17418-9" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1.96261,0,0,1.09426,-74.6625,-21.1211)" cx="77.5625" cy="152.51079" fx="77.5625" fy="152.51079" r="13.03125"/>
    <ns0:linearGradient id="linearGradient10599-4-0-8-1-6-9" ns1:collect="always">
      <ns0:stop id="stop10601-9-3-6-7-5-5-2" offset="0" style="stop-color: rgb(255, 255, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop10603-3-0-1-5-1-4" offset="1" style="stop-color: rgb(255, 255, 255); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:filter color-interpolation-filters="sRGB" id="filter10631-9-5-7-4-7-2" ns1:collect="always">
      <ns0:feGaussianBlur id="feGaussianBlur10633-6-0-3-5-7-96" stdDeviation="0.5906498" ns1:collect="always"/>
    </ns0:filter>
    <ns1:path-effect effect="spiro" id="path-effect30869" is_visible="true"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6996-2">
      <ns0:path id="path6998-8" d="m 290.13291,107.02249 c -0.52316,-1.95241 -2.52999,-3.11107 -4.4824,-2.58791 -0.96349,0.25817 -1.73966,0.87495 -2.20981,1.67092 l -0.0311,-0.0182 -33.7284,55.3598 c -0.10281,0.17003 -0.19825,0.34177 -0.28097,0.52259 l 0.008,0.0245 -0.28755,0.49803 0.0621,0.0359 c -0.28822,0.89781 -0.33736,1.8833 -0.0752,2.86186 0.72658,2.71169 3.51384,4.32089 6.22554,3.5943 1.43104,-0.38344 2.54552,-1.34541 3.18122,-2.56271 l 0.0311,0.0182 0.28402,-0.7076 31.0997,-56.23417 c 0.34119,-0.74663 0.43404,-1.62082 0.20495,-2.47567 z" style="color:#000000;fill:none;stroke:#000000;stroke-width:2;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0" ns2:nodetypes="csccccccccscccccc"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath7139-5">
      <ns0:path style="color:#000000;fill:none;stroke:#000000;stroke-width:2;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 257,136.25 c -2.48528,0 -4.5,2.01472 -4.5,4.5 0,1.22647 0.48552,2.34456 1.28125,3.15625 l -0.0312,0.0312 25.75,24.375 c 0.16907,0.17638 0.34266,0.34436 0.53125,0.5 l 0.0312,0 0.5,0.5 0.0625,-0.0625 c 0.97462,0.62799 2.12939,1 3.375,1 3.45178,0 6.25,-2.79822 6.25,-6.25 0,-1.82164 -0.78781,-3.45138 -2.03125,-4.59375 l 0.0312,-0.0312 -0.75,-0.5625 -27.625,-21.53125 C 259.09687,136.63839 258.08816,136.25 257,136.25 z" id="path7141-9" ns1:connector-curvature="0"/>
    </ns0:clipPath>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient7040-3-2" id="linearGradient23681" gradientUnits="userSpaceOnUse" gradientTransform="translate(0,-11)" x1="274.03629" y1="135.51024" x2="269.89642" y2="188.14354"/>
    <ns0:linearGradient id="linearGradient7040-3-2" ns1:collect="always">
      <ns0:stop id="stop7042-5-4" offset="0" style="stop-color:#d6d6d2;stop-opacity:1"/>
      <ns0:stop id="stop7044-4-1" offset="1" style="stop-color:#44443d;stop-opacity:1"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient3149-9" id="linearGradient6529" gradientUnits="userSpaceOnUse" x1="15.737708" y1="40.104774" x2="20.413162" y2="29.15625"/>
    <ns0:linearGradient id="linearGradient3149-9" ns1:collect="always">
      <ns0:stop id="stop3151-9" offset="0" style="stop-color:white;stop-opacity:1;"/>
      <ns0:stop id="stop3153-1" offset="1" style="stop-color:white;stop-opacity:0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient4724-9" id="radialGradient10861-2" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.3448276,0,20.043241)" cx="-648.922" cy="32.674965" fx="-648.922" fy="32.674965" r="5.126524"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient4724-9">
      <ns0:stop style="stop-color:#2e3436;stop-opacity:1" offset="0" id="stop4726-7"/>
      <ns0:stop style="stop-color:#000000;stop-opacity:1" offset="1" id="stop4728-3"/>
    </ns0:linearGradient>
    <ns1:path-effect effect="spiro" id="path-effect30843" is_visible="true"/>
    <ns0:filter color-interpolation-filters="sRGB" ns1:collect="always" id="filter52127" x="-0.057684805" width="1.1153696" y="-0.13389868" height="1.2677974">
      <ns0:feGaussianBlur ns1:collect="always" stdDeviation="0.86301877" id="feGaussianBlur52129"/>
    </ns0:filter>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath15654">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path15656" ns2:cx="180.375" ns2:cy="183.625" ns2:rx="20.875" ns2:ry="20.875" d="m 201.25,183.625 a 20.875,20.875 0 1 1 -41.75,0 20.875,20.875 0 1 1 41.75,0 z" transform="translate(253.75,41.5)"/>
    </ns0:clipPath>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient15503" id="radialGradient30641" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.7540107,0,53.856283)" cx="434.75894" cy="229.38165" fx="434.75894" fy="229.38165" r="11.6875"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient15503">
      <ns0:stop style="stop-color:#ffffff;stop-opacity:1" offset="0" id="stop15505"/>
      <ns0:stop style="stop-color:#ffffff;stop-opacity:0" offset="1" id="stop15507"/>
    </ns0:linearGradient>
    <ns0:radialGradient r="46.177555" fy="152.54469" fx="154.30887" cy="152.54469" cx="154.30887" gradientTransform="matrix(3.8062827,-4.3447397e-8,2.2199035e-8,1.944784,116.22821,273.72246)" gradientUnits="userSpaceOnUse" id="radialGradient25776" ns4:href="#linearGradient5467" ns1:collect="always"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient5467">
      <ns0:stop style="stop-color:#ffffff;stop-opacity:1;" offset="0" id="stop5469"/>
      <ns0:stop style="stop-color:#ffffff;stop-opacity:0.7173913" offset="1" id="stop5471"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient7040-3-2" id="linearGradient7395" gradientUnits="userSpaceOnUse" gradientTransform="translate(0,-11)" x1="274.03629" y1="135.51024" x2="269.89642" y2="188.14354"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient15503" id="radialGradient7468" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.7540107,0,53.856283)" cx="434.75894" cy="229.38165" fx="434.75894" fy="229.38165" r="11.6875"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient8346" id="linearGradient8358" gradientUnits="userSpaceOnUse" x1="383.12347" y1="405.51575" x2="383.12347" y2="387.5"/>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask8354">
      <ns0:rect style="color:#000000;fill:url(#linearGradient8358);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:0.24697506;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect8356" width="438" height="55" x="144" y="359"/>
    </ns0:mask>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-3-1-7" id="linearGradient14910-9" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient id="linearGradient5716-3-1-7">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-0-3-8"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-0-39-8"/>
    </ns0:linearGradient>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns0:metadata id="metadata1530">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="bg" ns2:insensitive="true">
    <ns0:rect style="fill:url(#GNOME);" id="background" width="864" height="487" x="-17" y="-9" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer3" ns1:label="thumb actual" style="opacity:0.4">
    <ns0:g transform="matrix(0.62961616,0,0,0.62961616,12.09573,7.9266974)" style="display:inline" ns1:export-ydpi="90" ns1:export-xdpi="90" ns1:export-filename="/home/jimmac/gfx/redhat/redhat-ux/Products/RHEL/RHEL7/video-jingles/tex/desktop.png" id="g8118">
      <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 79.06066,57.414214 1120.87864,0 0,51.485276 c 0,0 -4.0279,-10.606597 -11.0989,-10.96015 L 89,99 c -4.59619,-0.353553 -9.93934,5.5 -9.93934,5.5 z" id="path8120" ns1:connector-curvature="0" ns2:nodetypes="ccccccc"/>
      <ns0:g id="g8122" transform="translate(11,0)">
        <ns0:rect y="58.273582" x="69.273582" height="599.45282" width="1119.4529" id="rect8124" style="color:#000000;fill:none;stroke:#000000;stroke-width:3.54716229000000016;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" d="m 1188.199,108.766 c 0,-5.89806 -4.7813,-10.6794 -10.6794,-10.6794 l -1097.99931,0 c -5.89809,0 -10.6794,4.78134 -10.6794,10.6794" style="fill:none;stroke:#000000;stroke-width:2.37319922000000005px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" id="path8126"/>
        <ns0:text ns2:linespacing="125%" id="text8128" y="84.187378" x="83.374763" style="font-size:21.26189422999999934px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" xml:space="preserve"><ns0:tspan y="84.187378" x="83.374763" id="tspan8130" ns2:role="line">Aktiviteter</ns0:tspan></ns0:text>
        <ns0:text ns2:linespacing="125%" id="text8136" y="84.187378" x="628.8465" style="font-size:21.26189422999999934px;font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;text-align:center;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell Bold" xml:space="preserve"><ns0:tspan y="84.187378" x="628.8465" id="tspan8138" ns2:role="line">14:30</ns0:tspan></ns0:text>
      </ns0:g>
      <ns0:g ns1:label="view-grid" id="g7362" transform="matrix(4,0,0,4,12,-591)" style="display:inline">
        <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" id="rect7364" width="16" height="16" x="20" y="276" ns1:label="a"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="279" x="23.0623" height="2" width="2.0000002" id="rect13363" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13365" width="2.0000002" height="2" x="27.0623" y="279" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="279" x="31.0623" height="2" width="2.0000002" id="rect13367" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13369" width="2.0000002" height="2" x="23.0623" y="283.01562" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="283.01562" x="27.0623" height="2" width="2.0000002" id="rect13371" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13373" width="2.0000002" height="2" x="31.0623" y="283.01562" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="287" x="23.0623" height="2" width="2.0000002" id="rect13375" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13377" width="2.0000002" height="2" x="27.0623" y="287" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="287" x="31.0623" height="2" width="2.0000002" id="rect13379" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      </ns0:g>
      <ns0:rect ry="3.9916313" rx="3.97597" y="449.98785" x="93.987839" height="48.024311" width="58.024311" id="rect17308" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:5.97568892999999957;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:path style="fill:url(#radialGradient17454);fill-opacity:1;fill-rule:nonzero;stroke:url(#linearGradient17456);stroke-width:2;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" d="m 152.5802,231.92088 c 0,15.42134 -12.53696,27.92288 -27.99964,27.92288 -15.4641,0 -28.00032,-12.5017 -28.00032,-27.92288 0,-15.42062 12.53622,-27.92088 28.00032,-27.92088 15.46268,0 27.99964,12.50026 27.99964,27.92088 l 0,0 z" id="path8610-8" ns1:connector-curvature="0"/>
      <ns0:g id="g8612-2" style="fill:url(#radialGradient17368-69);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8614-5" style="fill:url(#radialGradient17366-7);fill-opacity:1">
          <ns0:path d="m 44.0713,20.7144 c 0,0.2627 0,0 0,0 l -0.5449,0.6172 c -0.334,-0.3936 -0.709,-0.7246 -1.0898,-1.0703 l -0.8359,0.123 -0.7637,-0.8633 0,1.0684 0.6543,0.4951 0.4355,0.4932 0.582,-0.6582 c 0.1465,0.2744 0.291,0.5488 0.4365,0.8232 l 0,0.8223 -0.6553,0.7402 -1.1992,0.8232 -0.9082,0.9063 -0.582,-0.6602 0.291,-0.7402 -0.5811,-0.6582 -0.9814,-2.0977 -0.8359,-0.9453 -0.2188,0.2461 0.3281,1.1934 0.6172,0.6992 c 0.3525,1.0176 0.7012,1.9902 1.1641,2.9629 0.7178,0 1.3945,-0.0762 2.1074,-0.166 l 0,0.5762 -0.8721,2.1392 -0.7998,0.9043 -0.6543,1.4004 c 0,0.7676 0,1.5352 0,2.3027 l 0.2188,0.9063 -0.3633,0.4102 -0.8008,0.4941 -0.8359,0.6992 0.6914,0.7813 -0.9453,0.8242 0.1816,0.5332 -1.418,1.6055 -0.9443,0 -0.7998,0.4941 -0.5098,0 0,-0.6582 -0.2168,-1.3184 c -0.2813,-0.8262 -0.5742,-1.6465 -0.8721,-2.4668 0,-0.6055 0.0361,-1.2051 0.0723,-1.8105 l 0.3643,-0.8223 -0.5098,-0.9883 0.0371,-1.3574 -0.6914,-0.7813 0.3457,-1.1309 -0.5625,-0.6382 -0.9824,0 -0.3271,-0.3701 -0.9814,0.6177 -0.3994,-0.4536 -0.9092,0.7817 c -0.6172,-0.6997 -1.2354,-1.3989 -1.8535,-2.0981 l -0.7266,-1.7285 0.6543,-0.9863 -0.3633,-0.4111 0.7988,-1.8936 c 0.6563,-0.8164 1.3418,-1.5996 2.0352,-2.3857 l 1.2363,-0.3291 1.3809,-0.1641 0.9453,0.2471 1.3447,1.3564 0.4727,-0.5342 0.6533,-0.082 1.2363,0.4111 0.9453,0 0.6543,-0.5762 0.291,-0.4111 -0.6553,-0.4111 -1.0908,-0.082 c -0.3027,-0.4199 -0.584,-0.8613 -0.9434,-1.2344 l -0.3643,0.1641 -0.1455,1.0703 -0.6543,-0.7402 -0.1445,-0.8242 -0.7266,-0.5742 -0.292,0 0.7275,0.8223 -0.291,0.7402 -0.5811,0.1641 0.3633,-0.7402 -0.6553,-0.3281 -0.5801,-0.6582 -1.0918,0.2461 -0.1445,0.3281 -0.6543,0.4121 -0.3633,0.9053 -0.9082,0.4521 -0.4004,-0.4521 -0.4355,0 0,-1.4814 0.9453,-0.4941 0.7266,0 -0.1465,-0.5752 -0.5801,-0.5762 0.9805,-0.2061 0.5449,-0.6162 0.4355,-0.7412 0.8008,0 -0.2188,-0.5752 0.5098,-0.3291 0,0.6582 1.0898,0.2461 1.0898,-0.9043 0.0732,-0.4121 0.9443,-0.6577 c -0.3418,0.0425 -0.6836,0.0737 -1.0176,0.1646 l 0,-0.7411 0.3633,-0.8228 -0.3633,0 -0.7984,0.7402 -0.2188,0.4116 0.2188,0.5767 -0.3643,0.9863 -0.5811,-0.3291 -0.5078,-0.5752 -0.8008,0.5752 -0.291,-1.3159 1.3809,-0.9048 0,-0.4941 0.873,-0.5757 1.3809,-0.3296 0.9453,0.3296 1.7441,0.3291 -0.4355,0.4932 -0.9453,0 0.9453,0.9873 0.7266,-0.8223 0.2207,-0.3618 c 0,0 2.7871,2.498 4.3799,5.2305 1.5928,2.7334 2.3408,5.9551 2.3408,6.6094 l 0,0 0,0 z" id="path8616-1" style="fill:url(#radialGradient17364);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8618-5" style="fill:url(#radialGradient17374-8);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8620-0" style="fill:url(#radialGradient17372-7);fill-opacity:1">
          <ns0:path d="m 26.0703,9.2363 -0.0732,0.4932 0.5098,0.3291 0.8711,-0.5757 -0.4355,-0.4937 -0.582,0.3296 -0.29,-0.0825" id="path8622-7" style="fill:url(#radialGradient17370);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8624-0" style="fill:url(#radialGradient17380-2);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8626-1" style="fill:url(#radialGradient17378-0);fill-opacity:1">
          <ns0:path d="m 26.8701,5.8633 -1.8906,-0.7407 -2.1797,0.2466 -2.6904,0.7402 -0.5088,0.4941 1.6719,1.1514 0,0.6582 -0.6543,0.6582 0.873,1.729 0.5801,-0.3301 0.7285,-1.1514 c 1.123,-0.3472 2.1299,-0.7407 3.1973,-1.2344 l 0.873,-2.2212" id="path8628-7" style="fill:url(#radialGradient17376);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8630-6" style="fill:url(#radialGradient17386-08);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8632-6" style="fill:url(#radialGradient17384-5);fill-opacity:1">
          <ns0:path d="m 28.833,12.7749 -0.291,-0.7412 -0.5098,0.165 0.1465,0.9043 0.6543,-0.3281" id="path8634-3" style="fill:url(#radialGradient17382);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8636-6" style="fill:url(#radialGradient17392-3);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8638-5" style="fill:url(#radialGradient17390-6);fill-opacity:1">
          <ns0:path d="m 29.123,12.6089 -0.1455,0.9883 0.7998,-0.165 0.5811,-0.5752 -0.5088,-0.4941 C 29.6787,11.9078 29.4824,11.483 29.2685,11.0465 l -0.4355,0 0,0.4932 0.29,0.3291 0,0.7402" id="path8640-6" style="fill:url(#radialGradient17388);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8648-9" style="fill:url(#radialGradient17398-2);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8650-6" style="fill:url(#radialGradient17396-0);fill-opacity:1">
          <ns0:path d="m 16.7656,9.5649 0.7266,0.4937 0.582,0 0,-0.5757 -0.7266,-0.3291 -0.582,0.4111" id="path8652-5" style="fill:url(#radialGradient17394);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8654-2" style="fill:url(#radialGradient17404-3);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8656-7" style="fill:url(#radialGradient17402-4);fill-opacity:1">
          <ns0:path d="m 14.876,8.9072 -0.3638,0.9048 0.7271,0 0.3638,-0.8228 C 15.9166,8.7675 16.2286,8.5444 16.5479,8.331 l 0.7271,0.2471 c 0.4844,0.3291 0.9688,0.6582 1.4536,0.9868 L 19.4561,8.9072 18.6558,8.5781 18.292,7.8374 16.9111,7.6728 16.8383,7.2612 16.184,7.4262 15.8936,8.002 15.5298,7.2613 l -0.145,0.3291 0.0728,0.8228 -0.5816,0.494" id="path8658-7" style="fill:url(#radialGradient17400);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8660-4" style="fill:url(#radialGradient17410-8);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8662-6" style="fill:url(#radialGradient17408-3);fill-opacity:1">
          <ns0:path d="M 17.4922,6.8496 17.856,6.521 18.5831,6.3564 c 0.498,-0.2422 0.998,-0.4053 1.5264,-0.5762 l -0.29,-0.4937 -0.9385,0.1348 -0.4434,0.4419 -0.731,0.106 -0.6499,0.3052 -0.3159,0.1528 -0.1929,0.2583 0.9443,0.1641" id="path8664-4" style="fill:url(#radialGradient17406);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8666-7" style="fill:url(#radialGradient17416-8);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,91.24312,201.37384)">
        <ns0:g id="g8668-3" style="fill:url(#radialGradient17414-5);fill-opacity:1">
          <ns0:path d="m 18.7285,14.6665 0.4365,-0.6582 -0.6548,-0.4932 0.2183,1.1514" id="path8670-2" style="fill:url(#radialGradient17412);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:path style="opacity:0.53513495000000000;fill:url(#radialGradient17418);fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter10631-9-5-7-4-7)" d="m 64.625,130 c -0.05592,0.48975 -0.09375,0.99536 -0.09375,1.5 0,7.1928 5.838446,13.03125 13.03125,13.03125 7.192801,0 13.031249,-5.83846 13.03125,-13.03125 0,-0.50479 -0.0378,-1.0101 -0.09375,-1.5 -0.753425,6.47773 -6.258685,11.53125 -12.9375,11.53125 -6.679033,0 -12.184356,-5.05322 -12.9375,-11.53125 z" transform="matrix(1.9727163,0,0,1.9727163,-28.36936,-27.23144)" id="path8734-7" ns1:connector-curvature="0"/>
      <ns0:path style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" d="m 152.5802,231.92088 c 0,15.42134 -12.53696,27.92288 -27.99964,27.92288 -15.4641,0 -28.00032,-12.5017 -28.00032,-27.92288 0,-15.42062 12.53622,-27.92088 28.00032,-27.92088 15.46268,0 27.99964,12.50026 27.99964,27.92088 l 0,0 z" id="path8610-4-7" ns1:connector-curvature="0"/>
      <ns0:path ns1:connector-curvature="0" id="path8676-0" d="m 124.26768,206.8372 -3,0.3125 -3.625,1 -0.6875,0.6875 2.25,1.5625 0,0.875 -0.875,0.9375 1.1875,2.3125 0.8125,-0.4375 0.9375,-1.5625 c 1.52724,-0.47204 2.92338,-1.0163 4.375,-1.6875 l 1.1875,-3 -2.5625,-1 z m -7,0.1874 -1.3125,0.1874 -0.625,0.625 -0.9375,0.125 -0.9375,0.4375 -0.375,0.1874 -0.3125,0.375 1.3125,0.1874 0.5,-0.4375 1,-0.1874 c 0.67726,-0.3293 1.3439,-0.58016 2.0625,-0.8125 l -0.375,-0.6875 z m -5.875,2.6875 -0.1874,0.4375 0.125,1.125 -0.8125,0.6875 -0.5,1.25 1,0 0.5,-1.125 c 0.42634,-0.3014 0.81578,-0.58488 1.25,-0.875 l 1,0.3125 c 0.65878,0.44742 1.3407,0.86576 2,1.3125 l 1,-0.875 -1.125,-0.4375 -0.5,-1 -1.875,-0.25 -0.0624,-0.5625 -0.9375,0.25 -0.375,0.75 -0.5,-1 z m -2.375,0.9375 -0.5,1.1875 c 0,0 -0.78744,0.1976 -1,0.25 -2.7146,2.50076 -8.22572,7.8712 -9.5,18.0625 0.0504,0.2363 0.9375,1.625 0.9375,1.625 l 2.0625,1.25 2.0625,0.5625 0.9375,1.0625 1.375,1.0625 0.75,-0.125 0.625,0.25 0,0.1874 -0.8125,2.125 -0.5625,0.875 0.1874,0.4375 -0.5,1.6875 1.75,3.25 1.8125,1.5625 0.8125,1.125 -0.125,2.375 0.5625,1.3125 -0.5625,2.5625 c 0,0 -0.0758,-0.008 0,0.25 0.0764,0.25762 3.17848,1.9585 3.375,1.8125 0.1958,-0.1488 0.375,-0.25 0.375,-0.25 l -0.1874,-0.5625 0.8125,-0.75 0.25,-0.8125 1.3125,-0.4375 1,-2.5 -0.3125,-0.625 0.6875,-1 1.5,-0.375 0.75,-1.75 -0.1874,-2.25 1.1875,-1.6875 0.1874,-1.6875 c -1.62298,-0.80458 -3.20164,-1.60914 -4.8125,-2.4375 l -0.8125,-1.5625 -1.4375,-0.375 -0.8125,-2.125 -2,0.25 -1.6875,-1.25 -1.75,1.5625 0,0.25 c -0.53854,-0.1554 -1.20798,-0.1428 -1.6875,-0.4375 l -0.375,-1.125 0,-1.25 -1.1875,0.125 c 0.099,-0.78338 0.1504,-1.59176 0.25,-2.375 l -0.6875,0 -0.6875,0.9375 -0.6875,0.3125 -1,-0.5625 -0.0624,-1.25 0.1874,-1.3125 1.5,-1.125 1.1875,0 0.1874,-0.6875 1.5,0.375 1.0625,1.3125 0.1874,-2.25 1.875,-1.5625 0.6875,-1.6875 1.375,-0.5625 0.8125,-1.0625 1.8125,-0.375 0.875,-1.3125 -2.6875,0 1.6875,-0.8125 1.1875,0 1.6875,-0.5625 0.1874,-0.6875 -0.625,-0.5 -0.6875,-0.25 0.25,-0.6875 -0.5,-1 -1.1875,0.4375 0.1874,-0.875 -1.375,-0.8125 -1.125,1.9375 0.125,0.6875 -1.125,0.4375 -0.6875,1.4375 -0.25,-1.3125 -1.875,-0.8125 -0.3125,-1 2.4375,-1.4375 1.125,-1.0625 0.0624,-1.1875 -0.5625,-0.375 -0.8125,-0.0624 z m 27.6875,0 -1.875,0.4375 -1.1875,0.75 0,0.6875 -1.875,1.25 0.4375,1.75 1.0625,-0.75 0.6875,0.75 0.8125,0.5 0.5,-1.375 -0.3125,-0.75 0.3125,-0.5625 1.0625,-1.0624 0.5,0 -0.5,1.125 0,1.0625 c 0.45424,-0.1236 0.91016,-0.1922 1.375,-0.25 l -1.25,0.875 -0.125,0.5625 -1.5,1.25 -1.4375,-0.3125 0,-0.9375 -0.6875,0.4375 0.25,0.8125 -1.0625,0 -0.3125,0.4375 -0.3125,0.5625 -0.6875,0.8125 -1.375,0.3125 0.8125,0.75 0.1874,0.8125 -1,0 -1.25,0.6875 0,2 0.5625,0 0.5625,0.625 1.25,-0.625 0.4375,-1.25 0.9375,-0.5625 0.1874,-0.4375 1.5,-0.3125 0.75,0.875 0.875,0.4375 -0.4375,1 0.75,-0.1874 0.4375,-1 -1,-1.125 0.375,0 1,0.75 0.1874,1.125 0.875,1 0.1874,-1.4375 0.5,-0.25 c 0.48876,0.50724 0.90084,1.11664 1.3125,1.6875 l 1.5,0.125 0.8754,0.5624 -0.375,0.5625 -0.9375,0.75 -1.25,0 -1.6875,-0.5 -0.875,0.0624 -0.6875,0.75 -1.8125,-1.875 -1.25,-0.3125 -1.9375,0.25 -1.625,0.4375 c -0.943,1.06874 -1.91998,2.14006 -2.8125,3.25 l -1.0625,2.5625 0.5,0.5625 -0.875,1.3125 0.9375,2.375 c 0.84058,0.9506 1.72312,1.92372 2.5625,2.875 l 1.1875,-1.125 0.5625,0.625 1.375,-0.8125 0.4375,0.5 1.3125,0 0.75,0.875 -0.4375,1.5 0.9375,1.0625 -0.0624,1.875 0.6875,1.3125 -0.5,1.125 c -0.0492,0.82306 -0.0624,1.6768 -0.0624,2.5 0.40512,1.11524 0.80494,2.18924 1.1875,3.3125 l 0.25,1.8125 0,0.875 0.6875,0 1.125,-0.625 1.25,0 1.9375,-2.1875 -0.25,-0.75 1.3125,-1.125 -0.9375,-1.0625 1.125,-0.9375 1.0625,-0.6875 0.5,-0.5625 -0.3125,-1.1875 0,-3.125 0.9375,-1.9375 1.0625,-1.25 1.1875,-2.875 0,-0.8125 c -0.5689,0.0716 -1.13126,0.1458 -1.6875,0.1874 l 1.125,-1.1875 1.625,-1.125 0.9375,-1 0,-1.125 c -0.1978,-0.37306 -0.4258,-0.75194 -0.625,-1.125 l -0.75,0.9375 -0.625,-0.6875 -0.875,-0.6875 0,-1.4375 1,1.1875 1.1875,-0.1874 c 0.51788,0.46998 0.98328,0.90238 1.4375,1.4375 l 0.75,-0.8125 c 0,-0.88956 -1.02136,-5.2838 -3.1875,-9 -2.16614,-3.71496 -5.9375,-7.125 -5.9375,-7.125 l -0.3125,0.5 -1,1.125 -1.25,-1.3125 1.25,0 0.625,-0.6875 -2.375,-0.4375 -1.3125,-0.4375 z m -5.125,6.6876 -0.6875,-0.6875 c -0.23242,-0.61874 -0.52162,-1.15656 -0.8125,-1.75 l -0.5625,0 0,0.625 0.375,0.5 0,1 -0.1874,1.3125 1.0625,-0.1874 0.8124,-0.8126 z m -4.625,-5.25 -0.8125,0.4375 -0.375,-0.125 -0.125,0.6875 0.6875,0.4375 1.1875,-0.75 -0.5625,-0.6875 z m -13.0625,0.1874 -0.8125,0.5625 1,0.6875 0.8125,0 0,-0.75 -1,-0.5 z m 15.1875,3.9375 -0.6875,0.25 0.1874,1.1875 0.9375,-0.4375 -0.4375,-1 z m -13.625,2 0.3125,1.5625 0.5625,-0.875 -0.875,-0.6875 z m 25.8125,8.75 1.125,1.3125 1.375,2.8125 0.75,0.875 -0.375,1.0625 0.75,0.8125 c -0.35104,0.024 -0.7015,0.0624 -1.0625,0.0624 -0.62952,-1.32244 -1.08312,-2.67904 -1.5625,-4.0625 l -0.875,-0.9375 -0.4375,-1.625 0.3125,-0.3125 z" style="fill:none;stroke:#000000;stroke-width:1;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;display:inline"/>
      <ns0:g style="display:inline" transform="matrix(2,0,0,2,-512.41982,-695.7253)" id="g8015-7">
        <ns0:path ns1:connector-curvature="0" d="m 316.42825,459.38669 -11.96834,11.62653 5.33417,0.0423 c 0,0 -2.18563,4.34708 -2.18563,4.34708 -0.67784,2.03351 2.63833,3.03097 3.14671,1.50584 0,0 1.97571,-4.36731 1.97571,-4.36731 l 3.71077,3.8688 -0.0134,-17.02323 z" id="path3480-8-9-9" ns2:nodetypes="cccssccc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#ffffff;stroke-width:3;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:path ns1:connector-curvature="0" d="m 316.42825,459.38669 -11.96834,11.62653 5.33417,0.0423 c 0,0 -2.18563,4.34708 -2.18563,4.34708 -0.67784,2.03351 2.63833,3.03097 3.14671,1.50584 0,0 1.97571,-4.36731 1.97571,-4.36731 l 3.71077,3.8688 -0.0134,-17.02323 z" id="path3480-8-5" ns2:nodetypes="cccssccc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#000000;stroke-width:0.99999994000000003;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      </ns0:g>
      <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:6;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 107.07098,284 -6.57078,6 -0.002,52 46,0 -0.002,-52 -6.57076,-6 -32.85386,0 z" id="rect2846-2-0-5" ns2:nodetypes="ccccccc"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccc" id="path4185-68-9-7-8" d="m 118.5,306 0,2 10,0 0,-2" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:round;stroke-opacity:1;display:inline;enable-background:new"/>
      <ns0:path ns2:nodetypes="ccccccc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-6-9" d="m 106.5,299.25 0,-3.25 34,0 0,5.5 m 0,12.5 -34,0 0,-7.25" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cccccc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-3-4-8" d="m 140.5,318 0,18 -34,0 m 0,-8.25 0,-9.75 23.375,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccc" id="path4185-68-9-7-5-7" d="m 118.5,328 0,2 10,0 0,-2" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:round;stroke-opacity:1;display:inline;enable-background:new"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-6-4-5" d="m 106.5,292 34,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccccccccccccc" id="rect2846-7-2-9-3-1-8-2" d="m 112.41664,364 c -2.81678,0 -5.26374,1.4564 -6.5716,3.62502 l -2.17838,5.01922 c -0.74014,1.22884 -1.16666,2.65724 -1.16666,4.18268 l 0,36.80772 c 0,4.6344 3.90252,8.36536 8.74996,8.36536 l 24.50006,0 c 4.84746,0 8.74998,-3.73096 8.74998,-8.36536 l 0,-36.80772 c 0,-1.52544 -0.4265,-2.95384 -1.16666,-4.18268 l -2.17836,-5.01922 C 139.84708,365.4564 137.40014,364 134.58334,364 l -22.1667,0 z" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:5.99999952000000025;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#000000;stroke:#000000;stroke-width:0.99999994000000003;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 123.50006,377.5 c -2.93596,0 -5.6175,0.99962 -7.76812,2.6729 l -1.33646,0 c -0.50904,0 -0.91882,0.4098 -0.91882,0.91882 l 0,1.33646 c -1.67328,2.15062 -2.6729,4.83218 -2.6729,7.76812 0,2.93594 0.99962,5.61748 2.6729,7.76812 l 0,1.33644 c 0,0.50902 0.40978,0.91882 0.91882,0.91882 l 1.33646,0 c 2.15062,1.67326 4.83216,2.6729 7.76812,2.6729 2.93594,0 5.61748,-0.99964 7.76812,-2.6729 l 1.33642,0 c 0.50904,0 0.91884,-0.4098 0.91884,-0.91882 l 0,-1.33644 c 1.67328,-2.15064 2.6729,-4.83218 2.6729,-7.76812 0,-2.93594 -0.99962,-5.6175 -2.6729,-7.76812 l 0,-1.33646 c 0,-0.50902 -0.4098,-0.91882 -0.91884,-0.91882 l -1.33642,0 C 129.11754,378.49962 126.436,377.5 123.50006,377.5 z" id="path3861-6-2-2-7-4-1-1" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 123.5,380.19628 c -5.52284,0 -9.99996,4.47716 -9.99996,10 0,5.52284 4.47712,10 9.99996,10 5.52286,0 10,-4.47716 10,-10 0,-5.52284 -4.47714,-10 -10,-10 z" id="path3861-6-4-8-5-2-0-1" ns2:nodetypes="csssc" ns1:connector-curvature="0"/>
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path3861-6-1-6-2-1-0-0" ns2:cx="143.75" ns2:cy="155.25" ns2:rx="63.25" ns2:ry="63.25" d="m 207,155.25 c 0,34.93201 -28.31799,63.25 -63.25,63.25 C 108.81799,218.5 80.5,190.18201 80.5,155.25 80.5,120.31799 108.81799,92 143.75,92 178.68201,92 207,120.31799 207,155.25 z" transform="matrix(0.06649192,0,0,0.06649192,113.9418,379.87338)"/>
      <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path3861-6-1-3-8-2-2" ns2:cx="143.75" ns2:cy="155.25" ns2:rx="63.25" ns2:ry="63.25" d="m 207,155.25 c 0,34.93201 -28.31799,63.25 -63.25,63.25 C 108.81799,218.5 80.5,190.18201 80.5,155.25 80.5,120.31799 108.81799,92 143.75,92 178.68201,92 207,120.31799 207,155.25 z" transform="matrix(-0.04273932,0,0,-0.04157418,129.64378,396.34832)"/>
      <ns0:path ns2:nodetypes="csssc" ns1:connector-curvature="0" id="path5385-7-4-7-8-0" d="m 130.28688,414.83107 c -1.09244,-0.91719 -1.78689,-2.29303 -1.78689,-3.83107 0,-2.76143 2.23858,-5 5.00001,-5 2.76143,0 5,2.23857 5,5 0,0.70532 -0.14604,1.37654 -0.40953,1.98505" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-miterlimit:4;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" id="path8330" d="m 104.5,462 5,4 -5,4" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1;display:inline"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path8332" d="m 112.67678,472 6,0" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1;display:inline"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 223.5196,96.0866 -131.99931,0 c -5.89809,0 -10.6794,4.78134 -10.6794,10.6794" style="fill:none;stroke:#000000;stroke-width:5;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path17186"/>
      <ns0:rect ry="24.20339" rx="24.20339" y="121.79661" x="488.77966" height="48.40678" width="290.44067" id="rect11062-3" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:path transform="matrix(2.6034636,0,0,2.6005055,-53.49059,-862.05263)" d="m 311,386.5 c 0,1.933 -1.567,3.5 -3.5,3.5 -1.933,0 -3.5,-1.567 -3.5,-3.5 0,-1.933 1.567,-3.5 3.5,-3.5 1.933,0 3.5,1.567 3.5,3.5 z" ns2:ry="3.5" ns2:rx="3.5" ns2:cy="386.5" ns2:cx="307.5" id="path27918" style="color:#000000;fill:none;stroke:#000000;stroke-width:1.55467153000000002;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      <ns0:path ns2:nodetypes="cc" id="path27941" d="m 754.16168,150.12192 8.09967,8.09046" style="color:#000000;fill:none;stroke:#000000;stroke-width:4.04523087000000015;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns1:connector-curvature="0"/>
      <ns0:rect style="opacity:0.70638272000000002;color:#000000;fill:none;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect1431" width="32.361851" height="32.361847" x="733.91248" y="129.89575"/>
      <ns0:path ns2:nodetypes="cssssc" ns1:connector-curvature="0" id="rect17188" d="m 79.70338,191.5 75.59324,0 c 6.76067,0 12.20338,5.44271 12.20338,12.20338 l 0,371.59324 c 0,6.76067 -5.44271,12.20338 -12.20338,12.20338 l -75.59324,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:rect ry="0" rx="0" y="457.49716" x="100.49716" height="32.005657" width="45.005657" id="rect17310" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.99434202999999999;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
    </ns0:g>
    <ns0:g id="g12195" transform="matrix(0.71005248,0,0,0.71005248,-2.038404,-249.63702)">
      <ns0:path style="fill:url(#radialGradient17454-5);fill-opacity:1;fill-rule:nonzero;stroke:url(#linearGradient17456-9);stroke-width:2;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" d="m 312.5802,564.28306 c 0,15.42134 -12.53696,27.92288 -27.99964,27.92288 -15.4641,0 -28.00032,-12.5017 -28.00032,-27.92288 0,-15.42062 12.53622,-27.92088 28.00032,-27.92088 15.46268,0 27.99964,12.50026 27.99964,27.92088 l 0,0 z" id="path8610-8-4" ns1:connector-curvature="0"/>
      <ns0:g id="g8612-2-3" style="fill:url(#radialGradient30900);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8614-5-6" style="fill:url(#radialGradient30898);fill-opacity:1">
          <ns0:path d="m 44.0713,20.7144 c 0,0.2627 0,0 0,0 l -0.5449,0.6172 c -0.334,-0.3936 -0.709,-0.7246 -1.0898,-1.0703 l -0.8359,0.123 -0.7637,-0.8633 0,1.0684 0.6543,0.4951 0.4355,0.4932 0.582,-0.6582 c 0.1465,0.2744 0.291,0.5488 0.4365,0.8232 l 0,0.8223 -0.6553,0.7402 -1.1992,0.8232 -0.9082,0.9063 -0.582,-0.6602 0.291,-0.7402 -0.5811,-0.6582 -0.9814,-2.0977 -0.8359,-0.9453 -0.2188,0.2461 0.3281,1.1934 0.6172,0.6992 c 0.3525,1.0176 0.7012,1.9902 1.1641,2.9629 0.7178,0 1.3945,-0.0762 2.1074,-0.166 l 0,0.5762 -0.8721,2.1392 -0.7998,0.9043 -0.6543,1.4004 c 0,0.7676 0,1.5352 0,2.3027 l 0.2188,0.9063 -0.3633,0.4102 -0.8008,0.4941 -0.8359,0.6992 0.6914,0.7813 -0.9453,0.8242 0.1816,0.5332 -1.418,1.6055 -0.9443,0 -0.7998,0.4941 -0.5098,0 0,-0.6582 -0.2168,-1.3184 c -0.2813,-0.8262 -0.5742,-1.6465 -0.8721,-2.4668 0,-0.6055 0.0361,-1.2051 0.0723,-1.8105 l 0.3643,-0.8223 -0.5098,-0.9883 0.0371,-1.3574 -0.6914,-0.7813 0.3457,-1.1309 -0.5625,-0.6382 -0.9824,0 -0.3271,-0.3701 -0.9814,0.6177 -0.3994,-0.4536 -0.9092,0.7817 c -0.6172,-0.6997 -1.2354,-1.3989 -1.8535,-2.0981 l -0.7266,-1.7285 0.6543,-0.9863 -0.3633,-0.4111 0.7988,-1.8936 c 0.6563,-0.8164 1.3418,-1.5996 2.0352,-2.3857 l 1.2363,-0.3291 1.3809,-0.1641 0.9453,0.2471 1.3447,1.3564 0.4727,-0.5342 0.6533,-0.082 1.2363,0.4111 0.9453,0 0.6543,-0.5762 0.291,-0.4111 -0.6553,-0.4111 -1.0908,-0.082 c -0.3027,-0.4199 -0.584,-0.8613 -0.9434,-1.2344 l -0.3643,0.1641 -0.1455,1.0703 -0.6543,-0.7402 -0.1445,-0.8242 -0.7266,-0.5742 -0.292,0 0.7275,0.8223 -0.291,0.7402 -0.5811,0.1641 0.3633,-0.7402 -0.6553,-0.3281 -0.5801,-0.6582 -1.0918,0.2461 -0.1445,0.3281 -0.6543,0.4121 -0.3633,0.9053 -0.9082,0.4521 -0.4004,-0.4521 -0.4355,0 0,-1.4814 0.9453,-0.4941 0.7266,0 -0.1465,-0.5752 -0.5801,-0.5762 0.9805,-0.2061 0.5449,-0.6162 0.4355,-0.7412 0.8008,0 -0.2188,-0.5752 0.5098,-0.3291 0,0.6582 1.0898,0.2461 1.0898,-0.9043 0.0732,-0.4121 0.9443,-0.6577 c -0.3418,0.0425 -0.6836,0.0737 -1.0176,0.1646 l 0,-0.7411 0.3633,-0.8228 -0.3633,0 -0.7984,0.7402 -0.2188,0.4116 0.2188,0.5767 -0.3643,0.9863 -0.5811,-0.3291 -0.5078,-0.5752 -0.8008,0.5752 -0.291,-1.3159 1.3809,-0.9048 0,-0.4941 0.873,-0.5757 1.3809,-0.3296 0.9453,0.3296 1.7441,0.3291 -0.4355,0.4932 -0.9453,0 0.9453,0.9873 0.7266,-0.8223 0.2207,-0.3618 c 0,0 2.7871,2.498 4.3799,5.2305 1.5928,2.7334 2.3408,5.9551 2.3408,6.6094 l 0,0 0,0 z" id="path8616-1-5" style="fill:url(#radialGradient17364-2);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8618-5-9" style="fill:url(#radialGradient30904);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8620-0-3" style="fill:url(#radialGradient30902);fill-opacity:1">
          <ns0:path d="m 26.0703,9.2363 -0.0732,0.4932 0.5098,0.3291 0.8711,-0.5757 -0.4355,-0.4937 -0.582,0.3296 -0.29,-0.0825" id="path8622-7-7" style="fill:url(#radialGradient17370-0);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8624-0-5" style="fill:url(#radialGradient30908);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8626-1-2" style="fill:url(#radialGradient30906);fill-opacity:1">
          <ns0:path d="m 26.8701,5.8633 -1.8906,-0.7407 -2.1797,0.2466 -2.6904,0.7402 -0.5088,0.4941 1.6719,1.1514 0,0.6582 -0.6543,0.6582 0.873,1.729 0.5801,-0.3301 0.7285,-1.1514 c 1.123,-0.3472 2.1299,-0.7407 3.1973,-1.2344 l 0.873,-2.2212" id="path8628-7-5" style="fill:url(#radialGradient17376-6);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8630-6-1" style="fill:url(#radialGradient30912);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8632-6-4" style="fill:url(#radialGradient30910);fill-opacity:1">
          <ns0:path d="m 28.833,12.7749 -0.291,-0.7412 -0.5098,0.165 0.1465,0.9043 0.6543,-0.3281" id="path8634-3-6" style="fill:url(#radialGradient17382-0);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8636-6-5" style="fill:url(#radialGradient30916);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8638-5-0" style="fill:url(#radialGradient30914);fill-opacity:1">
          <ns0:path d="m 29.123,12.6089 -0.1455,0.9883 0.7998,-0.165 0.5811,-0.5752 -0.5088,-0.4941 C 29.6787,11.9078 29.4824,11.483 29.2685,11.0465 l -0.4355,0 0,0.4932 0.29,0.3291 0,0.7402" id="path8640-6-8" style="fill:url(#radialGradient17388-62);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8648-9-4" style="fill:url(#radialGradient30920);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8650-6-6" style="fill:url(#radialGradient30918);fill-opacity:1">
          <ns0:path d="m 16.7656,9.5649 0.7266,0.4937 0.582,0 0,-0.5757 -0.7266,-0.3291 -0.582,0.4111" id="path8652-5-0" style="fill:url(#radialGradient17394-9);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8654-2-5" style="fill:url(#radialGradient30924);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8656-7-0" style="fill:url(#radialGradient30922);fill-opacity:1">
          <ns0:path d="m 14.876,8.9072 -0.3638,0.9048 0.7271,0 0.3638,-0.8228 C 15.9166,8.7675 16.2286,8.5444 16.5479,8.331 l 0.7271,0.2471 c 0.4844,0.3291 0.9688,0.6582 1.4536,0.9868 L 19.4561,8.9072 18.6558,8.5781 18.292,7.8374 16.9111,7.6728 16.8383,7.2612 16.184,7.4262 15.8936,8.002 15.5298,7.2613 l -0.145,0.3291 0.0728,0.8228 -0.5816,0.494" id="path8658-7-2" style="fill:url(#radialGradient17400-9);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8660-4-0" style="fill:url(#radialGradient30928);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8662-6-7" style="fill:url(#radialGradient30926);fill-opacity:1">
          <ns0:path d="M 17.4922,6.8496 17.856,6.521 18.5831,6.3564 c 0.498,-0.2422 0.998,-0.4053 1.5264,-0.5762 l -0.29,-0.4937 -0.9385,0.1348 -0.4434,0.4419 -0.731,0.106 -0.6499,0.3052 -0.3159,0.1528 -0.1929,0.2583 0.9443,0.1641" id="path8664-4-4" style="fill:url(#radialGradient17406-0);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g8666-7-1" style="fill:url(#radialGradient30932);fill-opacity:1;fill-rule:nonzero;stroke-miterlimit:4;display:inline" transform="matrix(1.3141735,0,0,1.3137808,251.24312,533.73602)">
        <ns0:g id="g8668-3-8" style="fill:url(#radialGradient30930);fill-opacity:1">
          <ns0:path d="m 18.7285,14.6665 0.4365,-0.6582 -0.6548,-0.4932 0.2183,1.1514" id="path8670-2-2" style="fill:url(#radialGradient17412-86);fill-opacity:1" ns1:connector-curvature="0"/>
        </ns0:g>
      </ns0:g>
      <ns0:path style="opacity:0.53513495;fill:url(#radialGradient17418-9);fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter10631-9-5-7-4-7-2)" d="m 64.625,130 c -0.05592,0.48975 -0.09375,0.99536 -0.09375,1.5 0,7.1928 5.838446,13.03125 13.03125,13.03125 7.192801,0 13.031249,-5.83846 13.03125,-13.03125 0,-0.50479 -0.0378,-1.0101 -0.09375,-1.5 -0.753425,6.47773 -6.258685,11.53125 -12.9375,11.53125 -6.679033,0 -12.184356,-5.05322 -12.9375,-11.53125 z" transform="matrix(1.9727163,0,0,1.9727163,131.63064,305.13074)" id="path8734-7-6" ns1:connector-curvature="0"/>
      <ns0:path style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" d="m 312.5802,564.28306 c 0,15.42134 -12.53696,27.92288 -27.99964,27.92288 -15.4641,0 -28.00032,-12.5017 -28.00032,-27.92288 0,-15.42062 12.53622,-27.92088 28.00032,-27.92088 15.46268,0 27.99964,12.50026 27.99964,27.92088 l 0,0 z" id="path8610-4-7-2" ns1:connector-curvature="0"/>
      <ns0:path ns1:connector-curvature="0" id="path8676-0-3" d="m 284.26768,539.19938 -3,0.3125 -3.625,1 -0.6875,0.6875 2.25,1.5625 0,0.875 -0.875,0.9375 1.1875,2.3125 0.8125,-0.4375 0.9375,-1.5625 c 1.52724,-0.47204 2.92338,-1.0163 4.375,-1.6875 l 1.1875,-3 -2.5625,-1 z m -7,0.1874 -1.3125,0.1874 -0.625,0.625 -0.9375,0.125 -0.9375,0.4375 -0.375,0.1874 -0.3125,0.375 1.3125,0.1874 0.5,-0.4375 1,-0.1874 c 0.67726,-0.3293 1.3439,-0.58016 2.0625,-0.8125 l -0.375,-0.6875 z m -5.875,2.6875 -0.1874,0.4375 0.125,1.125 -0.8125,0.6875 -0.5,1.25 1,0 0.5,-1.125 c 0.42634,-0.3014 0.81578,-0.58488 1.25,-0.875 l 1,0.3125 c 0.65878,0.44742 1.3407,0.86576 2,1.3125 l 1,-0.875 -1.125,-0.4375 -0.5,-1 -1.875,-0.25 -0.0624,-0.5625 -0.9375,0.25 -0.375,0.75 -0.5,-1 z m -2.375,0.9375 -0.5,1.1875 c 0,0 -0.78744,0.1976 -1,0.25 -2.7146,2.50076 -8.22572,7.8712 -9.5,18.0625 0.0504,0.2363 0.9375,1.625 0.9375,1.625 l 2.0625,1.25 2.0625,0.5625 0.9375,1.0625 1.375,1.0625 0.75,-0.125 0.625,0.25 0,0.1874 -0.8125,2.125 -0.5625,0.875 0.1874,0.4375 -0.5,1.6875 1.75,3.25 1.8125,1.5625 0.8125,1.125 -0.125,2.375 0.5625,1.3125 -0.5625,2.5625 c 0,0 -0.0758,-0.008 0,0.25 0.0764,0.25762 3.17848,1.9585 3.375,1.8125 0.1958,-0.1488 0.375,-0.25 0.375,-0.25 l -0.1874,-0.5625 0.8125,-0.75 0.25,-0.8125 1.3125,-0.4375 1,-2.5 -0.3125,-0.625 0.6875,-1 1.5,-0.375 0.75,-1.75 -0.1874,-2.25 1.1875,-1.6875 0.1874,-1.6875 c -1.62298,-0.80458 -3.20164,-1.60914 -4.8125,-2.4375 l -0.8125,-1.5625 -1.4375,-0.375 -0.8125,-2.125 -2,0.25 -1.6875,-1.25 -1.75,1.5625 0,0.25 c -0.53854,-0.1554 -1.20798,-0.1428 -1.6875,-0.4375 l -0.375,-1.125 0,-1.25 -1.1875,0.125 c 0.099,-0.78338 0.1504,-1.59176 0.25,-2.375 l -0.6875,0 -0.6875,0.9375 -0.6875,0.3125 -1,-0.5625 -0.0624,-1.25 0.1874,-1.3125 1.5,-1.125 1.1875,0 0.1874,-0.6875 1.5,0.375 1.0625,1.3125 0.1874,-2.25 1.875,-1.5625 0.6875,-1.6875 1.375,-0.5625 0.8125,-1.0625 1.8125,-0.375 0.875,-1.3125 -2.6875,0 1.6875,-0.8125 1.1875,0 1.6875,-0.5625 0.1874,-0.6875 -0.625,-0.5 -0.6875,-0.25 0.25,-0.6875 -0.5,-1 -1.1875,0.4375 0.1874,-0.875 -1.375,-0.8125 -1.125,1.9375 0.125,0.6875 -1.125,0.4375 -0.6875,1.4375 -0.25,-1.3125 -1.875,-0.8125 -0.3125,-1 2.4375,-1.4375 1.125,-1.0625 0.0624,-1.1875 -0.5625,-0.375 -0.8125,-0.0624 z m 27.6875,0 -1.875,0.4375 -1.1875,0.75 0,0.6875 -1.875,1.25 0.4375,1.75 1.0625,-0.75 0.6875,0.75 0.8125,0.5 0.5,-1.375 -0.3125,-0.75 0.3125,-0.5625 1.0625,-1.0624 0.5,0 -0.5,1.125 0,1.0625 c 0.45424,-0.1236 0.91016,-0.1922 1.375,-0.25 l -1.25,0.875 -0.125,0.5625 -1.5,1.25 -1.4375,-0.3125 0,-0.9375 -0.6875,0.4375 0.25,0.8125 -1.0625,0 -0.3125,0.4375 -0.3125,0.5625 -0.6875,0.8125 -1.375,0.3125 0.8125,0.75 0.1874,0.8125 -1,0 -1.25,0.6875 0,2 0.5625,0 0.5625,0.625 1.25,-0.625 0.4375,-1.25 0.9375,-0.5625 0.1874,-0.4375 1.5,-0.3125 0.75,0.875 0.875,0.4375 -0.4375,1 0.75,-0.1874 0.4375,-1 -1,-1.125 0.375,0 1,0.75 0.1874,1.125 0.875,1 0.1874,-1.4375 0.5,-0.25 c 0.48876,0.50724 0.90084,1.11664 1.3125,1.6875 l 1.5,0.125 0.8754,0.5624 -0.375,0.5625 -0.9375,0.75 -1.25,0 -1.6875,-0.5 -0.875,0.0624 -0.6875,0.75 -1.8125,-1.875 -1.25,-0.3125 -1.9375,0.25 -1.625,0.4375 c -0.943,1.06874 -1.91998,2.14006 -2.8125,3.25 l -1.0625,2.5625 0.5,0.5625 -0.875,1.3125 0.9375,2.375 c 0.84058,0.9506 1.72312,1.92372 2.5625,2.875 l 1.1875,-1.125 0.5625,0.625 1.375,-0.8125 0.4375,0.5 1.3125,0 0.75,0.875 -0.4375,1.5 0.9375,1.0625 -0.0624,1.875 0.6875,1.3125 -0.5,1.125 c -0.0492,0.82306 -0.0624,1.6768 -0.0624,2.5 0.40512,1.11524 0.80494,2.18924 1.1875,3.3125 l 0.25,1.8125 0,0.875 0.6875,0 1.125,-0.625 1.25,0 1.9375,-2.1875 -0.25,-0.75 1.3125,-1.125 -0.9375,-1.0625 1.125,-0.9375 1.0625,-0.6875 0.5,-0.5625 -0.3125,-1.1875 0,-3.125 0.9375,-1.9375 1.0625,-1.25 1.1875,-2.875 0,-0.8125 c -0.5689,0.0716 -1.13126,0.1458 -1.6875,0.1874 l 1.125,-1.1875 1.625,-1.125 0.9375,-1 0,-1.125 c -0.1978,-0.37306 -0.4258,-0.75194 -0.625,-1.125 l -0.75,0.9375 -0.625,-0.6875 -0.875,-0.6875 0,-1.4375 1,1.1875 1.1875,-0.1874 c 0.51788,0.46998 0.98328,0.90238 1.4375,1.4375 l 0.75,-0.8125 c 0,-0.88956 -1.02136,-5.2838 -3.1875,-9 -2.16614,-3.71496 -5.9375,-7.125 -5.9375,-7.125 l -0.3125,0.5 -1,1.125 -1.25,-1.3125 1.25,0 0.625,-0.6875 -2.375,-0.4375 -1.3125,-0.4375 z m -5.125,6.6876 -0.6875,-0.6875 c -0.23242,-0.61874 -0.52162,-1.15656 -0.8125,-1.75 l -0.5625,0 0,0.625 0.375,0.5 0,1 -0.1874,1.3125 1.0625,-0.1874 0.8124,-0.8126 z m -4.625,-5.25 -0.8125,0.4375 -0.375,-0.125 -0.125,0.6875 0.6875,0.4375 1.1875,-0.75 -0.5625,-0.6875 z m -13.0625,0.1874 -0.8125,0.5625 1,0.6875 0.8125,0 0,-0.75 -1,-0.5 z m 15.1875,3.9375 -0.6875,0.25 0.1874,1.1875 0.9375,-0.4375 -0.4375,-1 z m -13.625,2 0.3125,1.5625 0.5625,-0.875 -0.875,-0.6875 z m 25.8125,8.75 1.125,1.3125 1.375,2.8125 0.75,0.875 -0.375,1.0625 0.75,0.8125 c -0.35104,0.024 -0.7015,0.0624 -1.0625,0.0624 -0.62952,-1.32244 -1.08312,-2.67904 -1.5625,-4.0625 l -0.875,-0.9375 -0.4375,-1.625 0.3125,-0.3125 z" style="fill:none;stroke:#000000;stroke-width:1;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;display:inline"/>
      <ns0:g transform="matrix(2,0,0,2,-352.41982,-363.36312)" id="g8015-7-0" style="display:inline">
        <ns0:path ns1:connector-curvature="0" d="m 316.42825,459.38669 -11.96834,11.62653 5.33417,0.0423 c 0,0 -2.18563,4.34708 -2.18563,4.34708 -0.67784,2.03351 2.63833,3.03097 3.14671,1.50584 0,0 1.97571,-4.36731 1.97571,-4.36731 l 3.71077,3.8688 -0.0134,-17.02323 z" id="path3480-8-9-9-5" ns2:nodetypes="cccssccc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#ffffff;stroke-width:3;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:path ns1:connector-curvature="0" d="m 316.42825,459.38669 -11.96834,11.62653 5.33417,0.0423 c 0,0 -2.18563,4.34708 -2.18563,4.34708 -0.67784,2.03351 2.63833,3.03097 3.14671,1.50584 0,0 1.97571,-4.36731 1.97571,-4.36731 l 3.71077,3.8688 -0.0134,-17.02323 z" id="path3480-8-5-0" ns2:nodetypes="cccssccc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#000000;stroke-width:0.99999994;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g12187" transform="matrix(0.66014572,0,0,0.66014572,281.03226,-274.9988)" ns1:label="files">
      <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:6;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 267.07098,616.36218 -6.57078,6 -0.002,52 46,0 -0.002,-52 -6.57076,-6 -32.85386,0 z" id="rect2846-2-0-5-5" ns2:nodetypes="ccccccc"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccc" id="path4185-68-9-7-8-7" d="m 278.5,638.36218 0,2 10,0 0,-2" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:round;stroke-opacity:1;display:inline;enable-background:new"/>
      <ns0:path ns2:nodetypes="ccccccc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-6-9-5" d="m 266.5,631.61218 0,-3.25 34,0 0,5.5 m 0,12.5 -34,0 0,-7.25" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cccccc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-3-4-8-4" d="m 300.5,650.36218 0,18 -34,0 m 0,-8.25 0,-9.75 23.375,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns1:connector-curvature="0" ns2:nodetypes="cccc" id="path4185-68-9-7-5-7-2" d="m 278.5,660.36218 0,2 10,0 0,-2" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:round;stroke-opacity:1;display:inline;enable-background:new"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="rect2846-4-5-0-6-8-6-4-5-8" d="m 266.5,624.36218 34,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:g>
    <ns0:g id="g23668" transform="matrix(0.66014572,0,0,0.66014572,-60.978215,-221.36197)">
      <ns0:path transform="matrix(0.96153846,0,0,0.96153846,133.63462,24.821622)" d="m 442.5,560.86218 c 0,16.2924 -13.2076,29.5 -29.5,29.5 -16.2924,0 -29.5,-13.2076 -29.5,-29.5 0,-16.2924 13.2076,-29.5 29.5,-29.5 16.2924,0 29.5,13.2076 29.5,29.5 z" ns2:ry="29.5" ns2:rx="29.5" ns2:cy="560.86218" ns2:cx="413" id="path23368" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6.24000025;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      <ns0:g ns1:transform-center-y="34.344176" ns1:transform-center-x="10.791579" transform="matrix(0.31132618,-0.02705993,0.02705993,0.31132618,416.64896,523.26137)" id="g7279" style="display:inline;enable-background:new">
        <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 353.89029,162.43914 c -0.8148,0 -1.50438,0.49404 -1.81876,1.1916 -0.01,0.0203 -0.0127,0.0426 -0.0207,0.0626 l -29.75544,65.2389 0.0208,0.0206 c -0.10568,0.19141 -0.16726,0.41393 -0.16726,0.64802 0,0.73893 0.59899,1.33796 1.33791,1.33796 0.51126,0 0.94549,-0.28936 1.17075,-0.71078 l 0.0626,-0.10453 c 0.0143,-0.0341 0.0303,-0.0692 0.0421,-0.10453 l 30.75888,-64.40268 0.0421,-0.0421 c 0.0962,-0.14236 0.15163,-0.31565 0.20906,-0.48082 0.007,-0.0144 0.0159,-0.0275 0.0207,-0.0421 0.0622,-0.19398 0.10452,-0.39144 0.10452,-0.60625 0,-1.10833 -0.89849,-2.00688 -2.00693,-2.00688 z" id="path7250" ns1:connector-curvature="0" ns2:nodetypes="cccccsscccccccscc"/>
      </ns0:g>
      <ns0:g transform="matrix(0.3118804,0.01966854,-0.01966854,0.3118804,489.29329,510.78749)" ns1:transform-center-y="-21.161415" ns1:transform-center-x="-4.9738117" id="g7209" style="display:inline;enable-background:new">
        <ns0:g style="fill:#000000;fill-opacity:1;stroke:none" id="g6973" clip-path="url(#clipPath6996-2)" transform="translate(-110,0)">
          <ns0:path ns2:nodetypes="csccccccccscccccc" ns1:connector-curvature="0" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 290.13291,107.02249 c -0.52316,-1.95241 -2.52999,-3.11107 -4.4824,-2.58791 -0.96349,0.25817 -1.73966,0.87495 -2.20981,1.67092 l -0.0311,-0.0182 -33.7284,55.3598 c -0.10281,0.17003 -0.19825,0.34177 -0.28097,0.52259 l 0.008,0.0245 -0.28755,0.49803 0.0621,0.0359 c -0.28822,0.89781 -0.33736,1.8833 -0.0752,2.86186 0.72658,2.71169 3.51384,4.32089 6.22554,3.5943 1.43104,-0.38344 2.54552,-1.34541 3.18122,-2.56271 l 0.0311,0.0182 0.28402,-0.7076 31.0997,-56.23417 c 0.34119,-0.74663 0.43404,-1.62082 0.20495,-2.47567 z" id="path6946"/>
          <ns0:path id="path6971" d="m 290.13291,107.02249 c -0.52316,-1.95241 -2.52999,-3.11107 -4.4824,-2.58791 -0.96349,0.25817 -1.73966,0.87495 -2.20981,1.67092 l -0.0311,-0.0182 -33.7284,55.3598 c -0.10281,0.17003 -0.19825,0.34177 -0.28097,0.52259 l 0.008,0.0245 -0.28755,0.49803 0.0621,0.0359 c -0.28822,0.89781 -0.33736,1.8833 -0.0752,2.86186 0.72658,2.71169 3.51384,4.32089 6.22554,3.5943 1.43104,-0.38344 2.54552,-1.34541 3.18122,-2.56271 l 0.0311,0.0182 0.28402,-0.7076 31.0997,-56.23417 c 0.34119,-0.74663 0.43404,-1.62082 0.20495,-2.47567 z" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0" ns2:nodetypes="csccccccccscccccc"/>
        </ns0:g>
        <ns0:g id="g7116" clip-path="url(#clipPath7139-5)" transform="translate(-140,0)">
          <ns0:path ns1:connector-curvature="0" id="path6937" d="m 257,136.25 c -2.48528,0 -4.5,2.01472 -4.5,4.5 0,1.22647 0.48552,2.34456 1.28125,3.15625 l -0.0312,0.0312 25.75,24.375 c 0.16907,0.17638 0.34266,0.34436 0.53125,0.5 l 0.0312,0 0.5,0.5 0.0625,-0.0625 c 0.97462,0.62799 2.12939,1 3.375,1 3.45178,0 6.25,-2.79822 6.25,-6.25 0,-1.82164 -0.78781,-3.45138 -2.03125,-4.59375 l 0.0312,-0.0312 -0.75,-0.5625 -27.625,-21.53125 C 259.09687,136.63839 258.08816,136.25 257,136.25 z" style="color:#000000;fill:url(#linearGradient23681);fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
          <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 257,136.25 c -2.48528,0 -4.5,2.01472 -4.5,4.5 0,1.22647 0.48552,2.34456 1.28125,3.15625 l -0.0312,0.0312 25.75,24.375 c 0.16907,0.17638 0.34266,0.34436 0.53125,0.5 l 0.0312,0 0.5,0.5 0.0625,-0.0625 c 0.97462,0.62799 2.12939,1 3.375,1 3.45178,0 6.25,-2.79822 6.25,-6.25 0,-1.82164 -0.78781,-3.45138 -2.03125,-4.59375 l 0.0312,-0.0312 -0.75,-0.5625 -27.625,-21.53125 C 259.09687,136.63839 258.08816,136.25 257,136.25 z" id="path7114" ns1:connector-curvature="0"/>
        </ns0:g>
        <ns0:path transform="matrix(0.26022189,0,0,0.26022189,-0.6833974,-113.79205)" d="m 600,1068 c 0,24.3005 -19.69947,44 -44,44 -24.30053,0 -44,-19.6995 -44,-44 0,-24.3005 19.69947,-44 44,-44 24.30053,0 44,19.6995 44,44 z" ns2:ry="44" ns2:rx="44" ns2:cy="1068" ns2:cx="556" id="path6909" style="fill:#000000;fill-opacity:1;stroke:none;display:inline;enable-background:new" ns2:type="arc"/>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g30877" transform="matrix(0.66014572,0,0,0.66014572,63.314075,-222.89132)">
      <ns0:path ns1:connector-curvature="0" ns1:original-d="m 478.18096,537.76522 -18.73833,18.73833 14.84924,8.30851 18.03123,-5.83363 0,-6.36397 z" ns1:path-effect="#path-effect30869" id="path30867" d="m 478.18096,537.76522 -18.73833,18.73833 14.84924,8.30851 18.03123,-5.83363 0,-6.36397 -14.14214,-14.84924" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:10;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:g transform="matrix(3.7500031,0,0,3.7521005,-830.66729,-1500.7311)" ns1:label="inkscape" id="g13277" style="display:inline">
        <ns0:path ns1:connector-curvature="0" id="path13254" d="m 348.94707,543.0052 c -0.45398,0 -0.8959,0.16964 -1.24379,0.52861 l -6.18785,6.37443 c -0.34097,0.35183 -0.52184,0.81575 -0.52861,1.27489 -1e-4,0.007 0,0.0234 0,0.031 -6e-5,1.36608 3.65031,0.04 3.98012,1.71022 0.17851,0.90395 -1.99006,0.48981 -1.99006,1.39927 0,1.06688 3.06954,0.3332 3.94903,1.21269 0.36128,0.87948 -1.17511,0.73753 -0.90174,1.55474 0.5152,0.53164 1.67415,0.23016 1.89678,1.08832 0.25429,0.98026 1.91986,0.81115 2.89181,0.0931 0.5152,-0.53162 -0.79505,-0.77436 -0.27984,-1.30597 0.51519,-0.53163 3.05996,-0.4241 3.07838,-1.58584 -0.24319,-0.72981 -1.19805,-0.84765 -1.21272,-1.71021 -0.0512,-0.73049 0.78195,-0.51683 3.42043,-1.2438 1.05503,-0.49441 1.09237,-0.75739 1.08832,-1.2127 -8e-5,-0.009 0,-0.0214 0,-0.031 -0.006,-0.45914 -0.21875,-0.92306 -0.5597,-1.27489 l -6.15676,-6.37443 c -0.34788,-0.35901 -0.78981,-0.52861 -1.2438,-0.52861 z m 0.12437,1.33708 c 0.46755,0.004 1.74874,1.58409 2.89182,2.76743 0.32152,0.42998 -0.12437,0.87065 -0.12437,0.87065 l -2.3943,-1.30598 -1.05723,1.43037 -0.93282,-1.39928 -0.55972,2.17664 -1.64802,-0.99504 0.43533,-0.55969 2.58086,-2.64306 c 0.19795,-0.2011 0.34952,-0.3456 0.80845,-0.34204 z m 7.08961,9.57719 c -0.12574,-0.004 -0.25257,0.006 -0.34204,0.031 -0.16865,0.0486 -0.96755,0.077 -0.90174,0.68409 0.72383,0.3034 1.82743,0.54491 1.95897,-0.0621 0.0988,-0.4552 -0.3379,-0.63905 -0.71519,-0.65297 z m -12.34461,2.02114 c -0.0702,0.008 -0.11793,0.036 -0.18656,0.0621 -0.54894,0.20872 -0.91708,0.64774 -0.40424,0.83956 0.51291,0.1918 0.85636,-0.0109 1.30597,-0.24876 0.44967,-0.23797 0.43675,-0.28133 0.40424,-0.37313 -0.0623,0.0125 -0.47121,-0.24203 -0.90174,-0.27987 -0.0717,-0.006 -0.14746,-0.008 -0.21767,0 z" style="fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none"/>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g12179" transform="matrix(0.67009649,0,0,0.67009649,188.8159,-265.61639)">
      <ns0:path ns2:nodetypes="ccccccccccccc" id="rect2846-7-2-9-3-1-8-2-9" d="m 272.41664,696.36218 c -2.81678,0 -5.26374,1.4564 -6.5716,3.62502 l -2.17838,5.01922 c -0.74014,1.22884 -1.16666,2.65724 -1.16666,4.18268 l 0,36.80772 c 0,4.6344 3.90252,8.36536 8.74996,8.36536 l 24.50006,0 c 4.84746,0 8.74998,-3.73096 8.74998,-8.36536 l 0,-36.80772 c 0,-1.52544 -0.4265,-2.95384 -1.16666,-4.18268 l -2.17836,-5.01922 c -1.3079,-2.16862 -3.75484,-3.62502 -6.57164,-3.62502 l -22.1667,0 z" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:5.99999952;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#000000;stroke:#000000;stroke-width:0.99999994;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 283.50006,709.86218 c -2.93596,0 -5.6175,0.99962 -7.76812,2.6729 l -1.33646,0 c -0.50904,0 -0.91882,0.4098 -0.91882,0.91882 l 0,1.33646 c -1.67328,2.15062 -2.6729,4.83218 -2.6729,7.76812 0,2.93594 0.99962,5.61748 2.6729,7.76812 l 0,1.33644 c 0,0.50902 0.40978,0.91882 0.91882,0.91882 l 1.33646,0 c 2.15062,1.67326 4.83216,2.6729 7.76812,2.6729 2.93594,0 5.61748,-0.99964 7.76812,-2.6729 l 1.33642,0 c 0.50904,0 0.91884,-0.4098 0.91884,-0.91882 l 0,-1.33644 c 1.67328,-2.15064 2.6729,-4.83218 2.6729,-7.76812 0,-2.93594 -0.99962,-5.6175 -2.6729,-7.76812 l 0,-1.33646 c 0,-0.50902 -0.4098,-0.91882 -0.91884,-0.91882 l -1.33642,0 c -2.15064,-1.67328 -4.83218,-2.6729 -7.76812,-2.6729 z" id="path3861-6-2-2-7-4-1-1-5" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 283.5,712.55846 c -5.52284,0 -9.99996,4.47716 -9.99996,10 0,5.52284 4.47712,10 9.99996,10 5.52286,0 10,-4.47716 10,-10 0,-5.52284 -4.47714,-10 -10,-10 z" id="path3861-6-4-8-5-2-0-1-4" ns2:nodetypes="csssc" ns1:connector-curvature="0"/>
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path3861-6-1-6-2-1-0-0-7" ns2:cx="143.75" ns2:cy="155.25" ns2:rx="63.25" ns2:ry="63.25" d="m 207,155.25 c 0,34.93201 -28.31799,63.25 -63.25,63.25 C 108.81799,218.5 80.5,190.18201 80.5,155.25 80.5,120.31799 108.81799,92 143.75,92 178.68201,92 207,120.31799 207,155.25 z" transform="matrix(0.06649192,0,0,0.06649192,273.9418,712.23556)"/>
      <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path3861-6-1-3-8-2-2-0" ns2:cx="143.75" ns2:cy="155.25" ns2:rx="63.25" ns2:ry="63.25" d="m 207,155.25 c 0,34.93201 -28.31799,63.25 -63.25,63.25 C 108.81799,218.5 80.5,190.18201 80.5,155.25 80.5,120.31799 108.81799,92 143.75,92 178.68201,92 207,120.31799 207,155.25 z" transform="matrix(-0.04273932,0,0,-0.04157418,289.64378,728.7105)"/>
      <ns0:path ns2:nodetypes="csssc" ns1:connector-curvature="0" id="path5385-7-4-7-8-0-4" d="m 290.28688,747.19325 c -1.09244,-0.91719 -1.78689,-2.29303 -1.78689,-3.83107 0,-2.76143 2.23858,-5 5.00001,-5 2.76143,0 5,2.23857 5,5 0,0.70532 -0.14604,1.37654 -0.40953,1.98505" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-miterlimit:4;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:g>
    <ns0:g id="g12173" transform="matrix(0.67009649,0,0,0.67009649,99.756825,-250.48223)" ns1:label="terminal">
      <ns0:rect ry="3.9916313" rx="3.97597" y="782.35004" x="253.98784" height="48.024311" width="58.024311" id="rect17308-9" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:5.97599983;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" id="path8330-5" d="m 264.5,794.36218 5,4 -5,4" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1;display:inline"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path8332-7" d="m 272.67678,804.36218 6,0" style="fill:none;stroke:#000000;stroke-width:2px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1;display:inline"/>
      <ns0:rect ry="0" rx="0" y="789.85938" x="260.49716" height="32.005657" width="45.005657" id="rect17310-8" style="color:#000000;fill:none;stroke:#000000;stroke-width:0.99434203;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
    </ns0:g>
    <ns0:g transform="matrix(1.1285839,0,0,1.1285839,371.62792,-6.8220215)" id="g4134" ns1:label="charmap">
      <ns0:g transform="matrix(1.0897521,0,0,1.0897521,-13.6138,-62.807336)" id="g4466">
        <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3.24021435;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:block;overflow:visible;enable-background:new" d="m 80.818419,284.98677 20.363171,0 c 1.76269,0 3.18175,1.40646 3.18175,3.1535 l 0,21.4438 c 0,1.74703 -1.41906,3.1535 -3.18175,3.1535 l -20.363171,0 c -1.762692,0 -3.181749,-1.40647 -3.181749,-3.1535 l 0,-21.4438 c 0,-1.74704 1.419057,-3.1535 3.181749,-3.1535 z" id="rect2960-9-7-86-2-4-6-4-1" ns1:connector-curvature="0" ns2:nodetypes="sssssssss"/>
        <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.5;stroke-miterlimit:4;marker:none;visibility:visible;display:block;overflow:visible;enable-background:new" d="m 99.5,291.29857 c 0,-0.79576 -0.63183,-1.43639 -1.41667,-1.43639 l -14.16666,0 c -0.78484,0 -1.41667,0.64063 -1.41667,1.43639 l 0,2.15736 m 0,9.21875 0,1.83862 c 0,0.79575 0.63183,1.43638 1.41667,1.43638 l 14.16666,0 c 0.78484,0 1.41667,-0.64063 1.41667,-1.43638 l 0,-3.6146" id="rect3835-9-4-3-3-7-7-1" ns1:connector-curvature="0" ns2:nodetypes="cssccccsssc"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:0.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="M 80.56816,308.87484 83,305.36218" id="path4281-5" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:0.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="M 100.67308,307.8718 99,305.36218" id="path4281-3-5" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:0.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="M 81.35769,288.25064 83,290.36218" id="path4301-9" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:0.5;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="M 101.31875,287.38093 99,290.36218" id="path4303-0" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
        <ns0:g transform="translate(5.0000024,27.999999)" style="font-size:14.08609581px;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-align:start;line-height:125%;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;font-family:Cantarell;-inkscape-font-specification:Cantarell" id="text17029">
          <ns0:path ns1:connector-curvature="0" d="m 90.682976,265.21578 -2.507325,2.2256 0.549358,0.69022 2.591841,-2.16926 -0.633874,-0.74656 m -1.436782,4.73293 c 0.845165,0 1.352266,0.26763 1.549471,0.80291 0.08452,0.22537 0.126775,0.56344 0.126775,1.05645 l 0,0.0564 c -1.04237,0.0282 -1.887538,0.12677 -2.56367,0.2958 -0.887423,0.23947 -1.662159,0.88743 -1.662159,2.01432 0,1.09871 1.000114,1.85936 2.183345,1.85936 0.760648,0 1.450868,-0.28172 2.084742,-0.80291 l 0.25355,0.63388 0.859251,0 0,-4.40895 c 0,-1.1128 -0.225378,-1.6199 -0.943768,-2.09883 -0.380324,-0.25355 -0.971941,-0.38032 -1.760762,-0.38032 -0.788821,0 -1.549471,0.14086 -2.281947,0.42258 l 0,0.9156 c 0.577529,-0.19721 1.577643,-0.36624 2.155172,-0.36624 m -1.408609,4.08497 c 0,-0.16904 0.05634,-0.32398 0.154947,-0.49302 0.225377,-0.36624 0.605702,-0.59161 1.126887,-0.7043 0.281722,-0.0564 0.873339,-0.0986 1.803021,-0.12678 l 0,1.6199 c -0.408497,0.39441 -0.873339,0.64796 -1.422696,0.74657 -0.154947,0.0282 -0.309894,0.0423 -0.450755,0.0423 -0.169033,0 -0.338067,-0.0282 -0.464841,-0.0845 -0.394411,-0.18312 -0.746563,-0.52119 -0.746563,-1.00011" id="path17034"/>
        </ns0:g>
      </ns0:g>
      <ns0:g transform="translate(41,64)" id="g5463-5-4-0"/>
    </ns0:g>
    <ns0:g id="g20818" transform="matrix(0.6509069,0,0,0.6509069,2.3447072,-126.76724)">
      <ns0:g transform="matrix(3.3710655,0,0,3.3710655,-202.84919,-139.88211)" ns1:label="miro" id="g105356" style="fill:#000000;fill-opacity:1;stroke:none;display:inline">
        <ns0:path d="m 194,256 c -7.99181,0 -10.64868,8.72576 -11,9.375 3.27017,3.4245 6.33118,4.625 10,4.625 2.64737,0 4.51382,-2.00722 5.3125,-4 0.54877,-1.36923 0.73215,-3.11278 0.65625,-7 -0.99898,-2 -3.96978,-3 -4.96875,-3 z m -7,4 7.71875,0 c 0.56616,0 0.70232,0.0584 1.15625,0.1875 0.79339,0.34029 1.09163,1.07816 1.125,1.75 0.024,1.11117 -0.007,2.95106 0,4.0625 l -2,0 0,-1 0,-2.71875 L 195,262 c 0,-0.554 -0.44657,-1 -1,-1 -0.55344,0 -1,0.446 -1,1 l 0,0.28125 0,2.71875 c 0.002,0.34659 0.002,0.73212 0,1 l -2,0 0,-0.25 0,-3.75 c 0,-0.554 -0.446,-1 -1,-1 -0.554,0 -1,0.446 -1,1 -0.0181,0.50626 -0.006,1.25319 0,2 l 0,1 0,0.65625 0,0.0937 c 1.4e-4,0.0897 5e-4,0.18669 0,0.25 l -2,0 0,-6 z" ns1:href="#path17600" id="path20816" style="fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:3.5597055;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline;enable-background:new" ns4:href="#path17600" ns1:original="M 194 256 C 186.00819 256 183.35132 264.72576 183 265.375 C 186.27017 268.7995 189.33118 270 193 270 C 195.64737 270 197.51382 267.99278 198.3125 266 C 198.86127 264.63077 199.04465 262.88722 198.96875 259 C 197.96977 257 194.99897 256 194 256 z M 187 260 L 194.71875 260 C 195.28491 260 195.42107 260.0584 195.875 260.1875 C 196.66839 260.52779 196.96663 261.26566 197 261.9375 C 197.024 263.04867 196.993 264.88856 197 266 L 195 266 L 195 265 L 195 262.28125 L 195 262 C 195 261.446 194.55343 261 194 261 C 193.44656 261 193 261.446 193 262 L 193 262.28125 L 193 265 C 193.002 265.34659 193.002 265.73212 193 266 L 191 266 L 191 265.75 L 191 262 C 191 261.446 190.554 261 190 261 C 189.446 261 189 261.446 189 262 C 188.9819 262.50626 188.994 263.25319 189 264 L 189 265 L 189 265.65625 L 189 265.75 C 189.00014 265.8397 189.0005 265.93669 189 266 L 187 266 L 187 260 z " ns1:radius="0" ns2:type="inkscape:offset"/>
        <ns0:path ns1:connector-curvature="0" id="path17600" d="m 194.0002,256 c -7.99181,0 -10.64868,8.72576 -11,9.375 3.27017,3.4245 6.33118,4.625 10,4.625 2.64737,0 4.51382,-2.00722 5.3125,-4 0.54877,-1.36923 0.73215,-3.11278 0.65625,-7 -0.99898,-2 -3.96978,-3 -4.96875,-3 z m -7,4 7.71875,0 c 0.56616,0 0.70232,0.0584 1.15625,0.1875 0.79339,0.34029 1.09163,1.07816 1.125,1.75 0.024,1.11117 -0.007,2.95106 0,4.0625 l -2,0 0,-1 0,-2.71875 0,-0.28125 c 0,-0.554 -0.44657,-1 -1,-1 -0.55344,0 -1,0.446 -1,1 l 0,0.28125 0,2.71875 c 0.002,0.34659 0.002,0.73212 0,1 l -2,0 0,-0.25 0,-3.75 c 0,-0.554 -0.446,-1 -1,-1 -0.554,0 -1,0.446 -1,1 -0.0181,0.50626 -0.006,1.25319 0,2 l 0,1 0,0.65625 0,0.0937 c 1.4e-4,0.0897 5e-4,0.18669 0,0.25 l -2,0 0,-6 z" style="fill:#ffffff;fill-opacity:1;stroke:none;display:inline;enable-background:new"/>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g30613" transform="matrix(0.67009649,0,0,0.67009649,-91.638557,-211.64033)">
      <ns0:path d="m 415.5,624.875 c -3.80438,0 -6.875,0.82143 -6.875,1.84375 l 0,36.1875 c 0,1.02233 3.07062,1.84375 6.875,1.84375 l 39.4375,0 c 3.80437,0 6.875,-0.82142 6.875,-1.84375 l 0,-36.1875 c 0,-1.02232 -3.07063,-1.84375 -6.875,-1.84375 l -7.375,0 -0.0937,0.46875 -9.25,0.0312 -0.125,-0.5 -22.59375,0 z" ns1:href="#rect19224" id="path30591" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns4:href="#rect19224" ns1:original="M 415.5 624.875 C 411.69562 624.875 408.625 625.69643 408.625 626.71875 L 408.625 662.90625 C 408.625 663.92858 411.69562 664.75 415.5 664.75 L 454.9375 664.75 C 458.74187 664.75 461.8125 663.92858 461.8125 662.90625 L 461.8125 626.71875 C 461.8125 625.69643 458.74187 624.875 454.9375 624.875 L 447.5625 624.875 L 447.46875 625.34375 L 438.21875 625.375 L 438.09375 624.875 L 415.5 624.875 z " ns1:radius="0" ns2:type="inkscape:offset"/>
      <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:6;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 415.50021,624.86773 22.58279,0.008 0.13613,0.48403 9.24186,-0.0303 0.10588,-0.46134 7.38138,0 c 3.80437,0 6.8671,0.82302 6.8671,1.84534 l 0,36.18087 c 0,1.02233 -3.06273,1.84535 -6.8671,1.84535 l -39.44804,0 c -3.80438,0 -6.86711,-0.82302 -6.86711,-1.84535 l 0,-36.18087 c 0,-1.02232 3.06273,-1.84534 6.86711,-1.84534 z" id="rect19224" ns1:connector-curvature="0" ns2:nodetypes="sccccssssssss"/>
      <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:4.13201761;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter52127);enable-background:new" d="m 112.3125,52.53125 c -9.91951,0 -17.96875,2.850005 -17.96875,6.34375 0,1.933127 2.464014,3.652134 6.34375,4.8125 L 98.375,66.5 106,68 l 2.875,-2.53125 c 0.6345,0.02389 1.53499,0.21875 2.1875,0.21875 11.16951,0 19.1875,-3.318755 19.1875,-6.8125 0,-3.493745 -8.01799,-6.34375 -17.9375,-6.34375 z" transform="matrix(0.24201252,0,0,0.24201252,397.84496,613.66803)" id="path16978" ns1:connector-curvature="0" ns2:nodetypes="ssccccsss"/>
      <ns0:g transform="matrix(0.37915538,0,0,0.37915538,374.62159,591.25572)" id="g17331">
        <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.55063653;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter16757-8);enable-background:new" d="m 153.25,84.866387 42,0 1.6875,9.258613 -43.75,0 z" id="rect17096" ns1:connector-curvature="0" ns2:nodetypes="ccccc"/>
        <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.39318216;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter16757-8);enable-background:new" id="path17138" ns2:cx="182.6875" ns2:cy="87.5625" ns2:rx="3.4375" ns2:ry="1.5625" d="m 186.125,87.5625 c 0,0.862945 -1.53902,1.5625 -3.4375,1.5625 -1.89848,0 -3.4375,-0.699555 -3.4375,-1.5625 0,-0.862945 1.53902,-1.5625 3.4375,-1.5625 1.89848,0 3.4375,0.699555 3.4375,1.5625 z" transform="matrix(1.1740571,0,0,1.6705259,-40.505155,-57.027801)"/>
        <ns0:g clip-path="none" id="g17193" transform="matrix(-1,0,0.19314882,1,337.86402,0)">
          <ns0:path transform="matrix(1,0,0,0.92018529,0.25,7.5447954)" ns2:nodetypes="cscccsccc" ns1:connector-curvature="0" id="path17484" d="m 161.44607,93.616606 c 0,0 -0.78005,-0.459575 -0.73974,-0.90054 0.0572,-0.62659 -0.1991,-1.501402 1.21733,-1.474766 l 5.94382,-0.0055 -0.0833,-12.140633 -4.68188,-0.09685 c -3.45297,-0.07143 -3.18065,2.428014 -3.18065,2.428014 l -0.0623,12.190276 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.55063653;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" clip-path="none"/>
        </ns0:g>
        <ns0:g transform="translate(-6.10467,0)" id="g17494" clip-path="none">
          <ns0:path clip-path="none" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.55063653;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 161.44607,93.616606 c 0,0 -0.78005,-0.459575 -0.73974,-0.90054 0.0572,-0.62659 -0.1991,-1.501402 1.21733,-1.474766 l 5.94382,-0.0055 -0.0833,-12.140633 -4.68188,-0.09685 c -3.45297,-0.07143 -3.18065,2.428014 -3.18065,2.428014 l -0.0623,12.190276 z" id="path17496" ns1:connector-curvature="0" ns2:nodetypes="cscccsccc" transform="matrix(1,0,0,0.92018529,0,7.5447954)"/>
        </ns0:g>
      </ns0:g>
      <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:4.01754808;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path17064" ns2:cx="69.125" ns2:cy="83.5" ns2:rx="18.625" ns2:ry="6.5" d="M 87.75,83.5 C 87.75,87.089851 79.411303,90 69.125,90 58.838697,90 50.5,87.089851 50.5,83.5 50.5,79.910149 58.838697,77 69.125,77 79.411303,77 87.75,79.910149 87.75,83.5 z" transform="matrix(0.2742272,0,0,0.22592655,436.28476,607.87482)"/>
      <ns0:g transform="matrix(0.26269733,0,0,0.26269733,398.17699,601.56142)" id="g15942">
        <ns0:path transform="matrix(0.73543852,0,0,0.73543852,47.808877,47.521858)" d="m 199.25,179.625 c 0,11.80509 -9.56991,21.375 -21.375,21.375 -11.80509,0 -21.375,-9.56991 -21.375,-21.375 0,-11.80509 9.56991,-21.375 21.375,-21.375 11.80509,0 21.375,9.56991 21.375,21.375 z" ns2:ry="21.375" ns2:rx="21.375" ns2:cy="179.625" ns2:cx="177.875" id="path15830-8" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.23782039;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
        <ns0:g id="g15864" transform="matrix(0.70175439,0,0,0.70175439,53.274123,53.572369)"/>
        <ns0:g id="g15595" clip-path="url(#clipPath15654)" transform="matrix(1.2642868,0,0,1.2642868,-370.38728,-93.77475)">
          <ns0:g id="g15812" transform="translate(0,6)"/>
          <ns0:g id="g15702" transform="translate(0,-3)">
            <ns0:path transform="matrix(0.82352941,0,0,1,76.213235,4)" d="m 446.75,218.9375 c 0,4.86701 -5.23267,8.8125 -11.6875,8.8125 -6.45483,0 -11.6875,-3.94549 -11.6875,-8.8125 0,-4.86701 5.23267,-8.8125 11.6875,-8.8125 6.45483,0 11.6875,3.94549 11.6875,8.8125 z" ns2:ry="8.8125" ns2:rx="11.6875" ns2:cy="218.9375" ns2:cx="435.0625" id="path15698" style="color:#000000;fill:#191025;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
            <ns0:path transform="matrix(0.66251783,0,0,0.88269156,146.26334,26.183217)" d="m 446.75,218.9375 c 0,4.86701 -5.23267,8.8125 -11.6875,8.8125 -6.45483,0 -11.6875,-3.94549 -11.6875,-8.8125 0,-4.86701 5.23267,-8.8125 11.6875,-8.8125 6.45483,0 11.6875,3.94549 11.6875,8.8125 z" ns2:ry="8.8125" ns2:rx="11.6875" ns2:cy="218.9375" ns2:cx="435.0625" id="path15501" style="color:#000000;fill:url(#radialGradient30641);fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
            <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path15431" ns2:cx="434.5" ns2:cy="218.5" ns2:rx="5.5" ns2:ry="5.5" d="m 440,218.5 c 0,3.03757 -2.46243,5.5 -5.5,5.5 -3.03757,0 -5.5,-2.46243 -5.5,-5.5 0,-3.03757 2.46243,-5.5 5.5,-5.5 3.03757,0 5.5,2.46243 5.5,5.5 z" transform="matrix(1.1363636,0,0,1.1363636,-59.25,-31.545455)"/>
            <ns0:path id="path15427" d="m 424.58196,217.89188 c -0.007,-0.13515 -0.0168,-0.26536 -0.0168,-0.40215 0,-4.53716 4.34257,-8.77776 9.62229,-8.77776 5.27973,0 9.4973,4.2406 9.4973,8.77776 0,0.13679 -0.009,0.267 -0.0168,0.40215 -0.2474,-4.34766 -4.48503,-6.62561 -9.60557,-6.62561 -5.12056,0 -9.23319,2.27795 -9.48059,6.62561 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns1:connector-curvature="0" ns2:nodetypes="cssscscc"/>
            <ns0:g id="g15449" transform="matrix(0.8813906,0,0,0.8813906,53.848934,25.653047)">
              <ns0:path transform="matrix(1.1582075,-0.27647923,0,1.1582075,-91.614292,75.799371)" d="m 452.75,224.25 c 0,1.51878 -1.45507,2.75 -3.25,2.75 -1.79493,0 -3.25,-1.23122 -3.25,-2.75 0,-1.51878 1.45507,-2.75 3.25,-2.75 1.79493,0 3.25,1.23122 3.25,2.75 z" ns2:ry="2.75" ns2:rx="3.25" ns2:cy="224.25" ns2:cx="449.5" id="path15433" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
            </ns0:g>
          </ns0:g>
        </ns0:g>
      </ns0:g>
      <ns0:path transform="matrix(1.0487678,0,0,1.0487678,45.282304,-29.015526)" d="m 393,646.23718 c 0,6.48935 -5.26065,11.75 -11.75,11.75 -6.48935,0 -11.75,-5.26065 -11.75,-11.75 0,-6.48934 5.26065,-11.75 11.75,-11.75 6.48935,0 11.75,5.26066 11.75,11.75 z" ns2:ry="11.75" ns2:rx="11.75" ns2:cy="646.23718" ns2:cx="381.25" id="path30589" style="color:#000000;fill:#ffffff;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:9.07692337;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.55063653;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 415.82612,622.52874 c -0.0849,0 -0.16819,1.7e-4 -0.25212,10e-4 l -0.112,0.1216 -0.16808,-0.11356 c -0.17181,0.006 -0.33805,0.0152 -0.50424,0.0272 l -0.056,0.1247 -0.21477,-0.10242 c -0.16394,0.0151 -0.32406,0.0339 -0.48089,0.0543 l 0,0.1264 -0.26146,-0.0896 c -0.15497,0.0238 -0.30674,0.0495 -0.45288,0.0784 l 0.0607,0.1247 -0.2988,-0.0752 c -0.14157,0.0317 -0.27973,0.066 -0.41087,0.10242 l 0.1168,0.1199 -0.32683,-0.0576 c -0.12555,0.0389 -0.24603,0.0801 -0.3595,0.12315 l 0.16808,0.11201 -0.35017,-0.0399 c -0.10608,0.0449 -0.20619,0.0923 -0.2988,0.14078 l 0.21943,0.10242 -0.36418,-0.0209 c -0.0843,0.0501 -0.15924,0.10213 -0.22877,0.15514 l 0.26146,0.0896 -0.36884,0 c -0.06,0.0538 -0.11454,0.10862 -0.15875,0.16474 l 0.29881,0.0736 -0.36416,0.0192 c -0.035,0.057 -0.0614,0.11384 -0.0794,0.17275 l 0.3315,0.0575 -0.35485,0.0384 c -0.004,0.0288 -0.004,0.0573 -0.004,0.0863 0,0.0291 5.2e-4,0.0575 0.004,0.0863 l 0.35485,0.0384 -0.3315,0.0575 c 0.0181,0.0588 0.0444,0.11581 0.0794,0.17273 l 0.36416,0.0192 -0.29881,0.0735 c 0.0443,0.0561 0.0987,0.11102 0.15875,0.16475 l 0.36884,0 -0.26146,0.0896 c 0.0695,0.053 0.14446,0.10509 0.22877,0.15514 l 0.36418,-0.0207 -0.21943,0.10241 c 0.0925,0.0485 0.19275,0.0958 0.2988,0.14078 l 0.35017,-0.0399 -0.16808,0.112 c 0.11342,0.043 0.234,0.0843 0.3595,0.12315 l 0.32683,-0.0576 -0.1168,0.11991 c 0.13118,0.0364 0.2693,0.0707 0.41087,0.10241 l 0.2988,-0.0752 -0.0607,0.1247 c 0.14614,0.0289 0.29791,0.0546 0.45288,0.0784 l 0.26146,-0.0896 0,0.12639 c 0.15683,0.0206 0.31695,0.0392 0.48089,0.0543 l 0.21477,-0.10241 0.056,0.12469 c 0.16619,0.0127 0.33243,0.021 0.50424,0.0272 l 0.16808,-0.11356 0.112,0.1216 c 0.0839,10e-4 0.16716,10e-4 0.25212,10e-4 0.0849,0 0.16819,-1.1e-4 0.25212,-10e-4 l 0.112,-0.1216 0.16808,0.11356 c 0.1718,-0.006 0.33805,-0.0152 0.50424,-0.0272 l 0.056,-0.12469 0.21477,0.10241 c 0.16394,-0.0151 0.32406,-0.0339 0.48089,-0.0543 l 0,-0.12639 0.26146,0.0896 c 0.15497,-0.0238 0.30673,-0.0495 0.45288,-0.0784 l -0.0607,-0.1247 0.29881,0.0752 c 0.14157,-0.0317 0.27972,-0.066 0.41086,-0.10241 l -0.11666,-0.11991 0.32682,0.0576 c 0.12554,-0.0389 0.24602,-0.0801 0.35951,-0.12315 l -0.16808,-0.112 0.35016,0.0399 c 0.10608,-0.0449 0.20619,-0.0923 0.29881,-0.14078 l -0.21943,-0.10241 0.36416,0.0207 c 0.0844,-0.0501 0.15926,-0.10199 0.22878,-0.15514 l -0.26146,-0.0896 0.36885,0 c 0.06,-0.0538 0.11454,-0.10862 0.15873,-0.16475 l -0.29881,-0.0735 0.36418,-0.0192 c 0.035,-0.057 0.0612,-0.11383 0.0794,-0.17273 l -0.3315,-0.0575 0.35485,-0.0384 c 0.004,-0.0288 0.004,-0.0573 0.004,-0.0863 0,-0.0291 -5.2e-4,-0.0575 -0.004,-0.0863 l -0.35485,-0.0384 0.3315,-0.0575 c -0.0181,-0.0588 -0.0444,-0.11581 -0.0794,-0.17275 l -0.36418,-0.0192 0.29881,-0.0736 c -0.0443,-0.0562 -0.0987,-0.11102 -0.15873,-0.16474 l -0.36885,0 0.26146,-0.0896 c -0.0695,-0.053 -0.14445,-0.10509 -0.22878,-0.15514 l -0.36416,0.0207 0.21943,-0.10241 c -0.0927,-0.0485 -0.19275,-0.0958 -0.29881,-0.14078 l -0.35016,0.0399 0.16808,-0.112 c -0.11356,-0.043 -0.23401,-0.0844 -0.35951,-0.12315 l -0.32682,0.0576 0.11666,-0.11991 c -0.13119,-0.0364 -0.26929,-0.0707 -0.41086,-0.10241 l -0.29881,0.0752 0.0607,-0.1247 c -0.14615,-0.0289 -0.29791,-0.0546 -0.45288,-0.0784 l -0.26146,0.0896 0,-0.12639 c -0.15683,-0.0206 -0.31695,-0.0392 -0.48089,-0.0543 l -0.21477,0.10241 -0.056,-0.12469 c -0.16619,-0.0127 -0.33244,-0.021 -0.50424,-0.0272 l -0.16808,0.11356 -0.112,-0.1216 c -0.0839,-0.001 -0.16714,-0.001 -0.25212,-0.001 z" id="path16671" ns1:connector-curvature="0"/>
      <ns0:path transform="matrix(-1,0,0,1,834.625,0)" ns2:open="true" ns2:end="7.609003" ns2:start="3.1415927" d="m 414.75,636.92468 c 0,-1.41523 1.14727,-2.5625 2.5625,-2.5625 1.41523,0 2.5625,1.14727 2.5625,2.5625 0,1.17585 -0.80026,2.20081 -1.941,2.48599" ns2:ry="2.5625" ns2:rx="2.5625" ns2:cy="636.92468" ns2:cx="417.3125" id="path30611" style="color:#000000;fill:#ffffff;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
    </ns0:g>
    <ns0:g style="display:inline" id="g68309" transform="matrix(0.73812401,0,0,0.73812401,450.6586,203.09701)" ns1:label="help">
      <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="cszsc" id="path3751" d="m 14.883007,5.3804864 c 0,4.5113247 -6.1837857,12.1788466 -7.884289,8.1726886 C 3.7280353,5.8478818 -1.1480278,12.785825 -3.4540023,8.2192786 -5.7318686,3.7083956 5.0017747,3.4589032 6.0524539,-0.76449404 7.5657882,-6.8476209 14.883007,0.86916191 14.883007,5.3804864 z" ns1:connector-curvature="0"/>
      <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="csszz" id="path3753" d="m 49.570335,7.2077552 c 5.552326,3.1568318 -4.054237,6.3454198 -8.406364,6.3454198 -4.352128,0 -7.88429,-3.6613639 -7.88429,-8.1726886 0,-4.51132449 6.299344,-8.4568909 10.364154,-5.69282488 4.004574,2.72310568 0.30796,4.32561458 5.9265,7.52009368 z" ns1:connector-curvature="0"/>
      <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="czzsc" id="path3755" d="M 14.883007,40.795492 C 10.153865,42.297569 9.5817611,52.389019 5.8507498,49.598133 1.9051658,46.646743 6.5683818,41.370391 0.39546008,42.207355 -5.749129,43.040477 -1.6161417,34.542357 6.998718,32.622802 c 4.247952,-0.946524 7.884289,3.661364 7.884289,8.17269 z" ns1:connector-curvature="0"/>
      <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="czzsz" id="path3757" d="m 48.695879,41.523268 c -6.690955,1.878845 -1.74186,7.467642 -6.494845,8.101936 -4.565071,0.60922 -6.451929,-4.759667 -7.063008,-8.829712 -0.607512,-4.046283 2.723221,-11.00695 6.025945,-8.17269 2.842221,2.439078 14.270309,7.008298 7.531908,8.900466 z" ns1:connector-curvature="0"/>
      <ns0:path style="fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:5.44904566;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" id="path1871" d="m 24.038299,-1.8893343 c -13.331156,0 -24.15066551,11.215268 -24.15066551,25.0340843 0,13.818818 10.81950951,25.034086 24.15066551,25.034086 13.331155,0 24.150665,-11.215268 24.150665,-25.034086 0,-13.8188163 -10.81951,-25.0340843 -24.150665,-25.0340843 z m 0,13.1758353 c 6.314752,-2e-6 11.439789,5.312505 11.439789,11.858249 0,6.545744 -5.125037,11.85825 -11.439789,11.85825 -6.314753,0 -11.439789,-5.312506 -11.439789,-11.85825 0,-6.545744 5.125036,-11.858249 11.439789,-11.858249 z" ns1:connector-curvature="0"/>
      <ns0:path ns2:nodetypes="ssssssssss" ns1:connector-curvature="0" d="m 24.038299,0.64151822 c -11.983426,0 -21.7091234,10.08144678 -21.7091234,22.50323178 0,12.421787 9.7256974,22.503233 21.7091234,22.503233 11.983425,0 21.709123,-10.081446 21.709123,-22.503233 0,-12.421785 -9.725698,-22.50323178 -21.709123,-22.50323178 z m 0,11.75499178 c 5.72365,-10e-7 10.368951,4.81522 10.368951,10.74824 0,5.93302 -4.645301,10.748241 -10.368951,10.748241 -5.723651,0 -10.368951,-4.815221 -10.368951,-10.748241 0,-5.93302 4.6453,-10.74824 10.368951,-10.74824 z" id="path68307" style="fill:#ffffff;fill-opacity:1;stroke:none"/>
      <ns0:path id="path2764" d="M 15.285859,2.4743562 C 10.300148,4.7510891 6.2906124,8.8924864 4.0942149,14.060578 c 4.5852109,-0.05424 7.5641511,2.312337 10.4742311,4.770797 1.039847,-2.439378 2.955558,-4.410322 5.308857,-5.488211 C 19.04958,9.2220694 17.608406,5.5277226 15.285859,2.4743562 z m 17.504879,0 c -2.236928,2.9126777 -4.141872,6.1687757 -4.591443,10.8688078 2.353298,1.077889 4.269009,3.048833 5.308856,5.488211 3.649601,-3.010131 7.184393,-4.998491 10.474231,-4.770797 C 41.785985,8.8924864 37.776449,4.7510891 32.790738,2.4743562 z M 14.568446,27.440332 c -3.491414,0.891924 -6.9828169,1.139291 -10.4742311,4.770797 2.1963975,5.16809 6.2059331,9.345358 11.1916441,11.622092 0.6226,-4.22438 1.814986,-8.080331 4.591444,-10.868809 -2.353299,-1.077889 -4.26901,-3.084703 -5.308857,-5.52408 z m 18.939705,0 c -1.039847,2.439377 -2.955558,4.446191 -5.308856,5.52408 2.320332,2.829279 3.711757,6.598889 4.591443,10.868809 4.985711,-2.276734 8.995247,-6.454002 11.191644,-11.622092 -2.4835,-2.795962 -6.191952,-4.133379 -10.474231,-4.770797 z" style="fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:g id="g30861" transform="matrix(0.67009649,0,0,0.67009649,131.3373,-275.87328)">
      <ns0:path d="m 388.37841,950.53882 c 0,6.9318 -5.57977,12.55114 -12.46276,12.55114 -6.88299,0 -12.46276,-5.61934 -12.46276,-12.55114 0,-6.93181 5.57977,-12.55115 12.46276,-12.55115 6.88299,0 12.46276,5.61934 12.46276,12.55115 z" ns2:ry="12.551146" ns2:rx="12.462757" ns2:cy="950.53882" ns2:cx="375.91565" id="path30859" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:12;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      <ns0:g transform="matrix(3.75,0,0,3.75,-789.66632,-1118.5571)" ns1:label="blender" id="g12660" style="display:inline">
        <ns0:path ns2:nodetypes="csccccsssccsccssccccsssss" style="fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:0.5333333;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 67.8125,328.0625 c -0.24052,0.0404 -0.472023,0.15754 -0.625,0.375 -0.305953,0.43491 -0.212493,1.03265 0.21875,1.34375 l 1.6875,1.21875 -1.28125,0 -1.0625,0 -3.71875,0 C 62.473823,331 62,331.44257 62,332 c 0,0.55743 0.473823,1 1.03125,1 l 2.903109,0 -4.432138,5.08839 c -0.419418,0.48332 -0.638516,1.14294 -0.189721,1.59911 0.448795,0.45617 1.143082,0.45207 1.5625,-0.0312 l 2.4375,-2.8125 c 0.510062,1.36413 1.653338,2.50504 3.21875,2.96875 2.640781,0.78227 5.458668,-0.61365 6.28125,-3.125 0.62887,-1.91995 -0.09979,-3.93258 -1.65625,-5.125 l -4.625,-3.34375 c -0.215622,-0.15555 -0.47823,-0.19664 -0.71875,-0.15625 z m 2.1875,4 c 1.656494,0 3,1.30442 3,2.9375 0,1.63308 -1.343506,2.96875 -3,2.96875 -1.656494,0 -3,-1.33567 -3,-2.96875 0,-1.63308 1.343506,-2.9375 3,-2.9375 z" transform="translate(241.0002,217)" id="rect12618" ns1:connector-curvature="0"/>
        <ns0:path ns2:type="arc" style="fill:#000000;fill-opacity:1;stroke:none" id="path12638" ns2:cx="69.09375" ns2:cy="333.98828" ns2:rx="0.9296875" ns2:ry="0.94140625" d="m 70.023437,333.98828 c 0,0.51993 -0.416235,0.94141 -0.929687,0.94141 -0.513452,0 -0.929688,-0.42148 -0.929688,-0.94141 0,-0.51992 0.416236,-0.94141 0.929688,-0.94141 0.513452,0 0.929687,0.42149 0.929687,0.94141 z" transform="matrix(1.8621708,0,0,1.7996949,182.32089,-49.374842)"/>
      </ns0:g>
    </ns0:g>
    <ns0:g id="g30890" transform="matrix(0.67009649,0,0,0.67009649,-20.649291,-204.63712)">
      <ns0:path id="path30882" d="m 461.875,611.625 c -12.70255,0 -23,10.29745 -23,23 0,12.70255 10.29745,23 23,23 2.01923,0 3.97777,-0.26129 5.84375,-0.75 -0.2175,-1.28287 -0.34375,-2.5927 -0.34375,-3.9375 0,-10.74315 7.23535,-19.82498 17.09375,-22.59375 C 482.45828,619.69241 473.11074,611.625 461.875,611.625 z m 0,17.25 c 3.17564,0 5.75,2.57436 5.75,5.75 0,3.17564 -2.57436,5.75 -5.75,5.75 -3.17564,0 -5.75,-2.57436 -5.75,-5.75 0,-3.17564 2.57436,-5.75 5.75,-5.75 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:10;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns1:connector-curvature="0"/>
      <ns0:g transform="matrix(3.75,0,0,3.75,-704.25078,-201.88856)" ns1:label="sound-juicer" id="g14313" style="display:inline">
        <ns0:rect style="fill:none;stroke:none" id="rect19048" width="16" height="16" x="303.00021" y="215"/>
        <ns0:path ns1:connector-curvature="0" id="path12550" d="m 310.96895,216 c -3.84231,0 -6.96875,3.18947 -6.96875,7.09375 0,3.90429 3.12644,6.9375 6.96875,6.9375 0.69879,0 1.35969,-0.11302 2,-0.3125 -0.41187,-1.9375 -0.42338,-3.03961 0.5,-4.71875 0.54324,-0.98785 1.74686,-2.96274 4.34375,-3.1875 C 317.31004,218.3938 314.46624,216 310.96895,216 z m 0.53125,1.0625 c 0.28659,0.0176 0.55406,0.11017 0.875,0.28125 0.66438,0.35416 0.99368,0.7203 0.8125,1.0625 l -1.03125,1.9375 c 0.95271,0.49213 1.625,1.48092 1.625,2.65625 0,1.65685 -1.3141,3 -2.90625,3 -0.25821,0 -0.51212,-0.0266 -0.75,-0.0937 l -0.5625,2.0625 c -0.11659,0.4319 -0.40529,0.55923 -1.15625,0.3125 -0.82913,-0.27249 -1.16906,-0.49422 -1.53125,-1.125 -0.37491,-0.65292 -0.46027,-1.14999 -0.125,-1.34375 l 1.8125,-1.03125 c -0.12379,-0.17416 -0.22663,-0.36296 -0.3125,-0.5625 l -1.84375,0.875 c -0.40383,0.19136 -0.66905,0.0752 -0.96875,-0.65625 -0.33084,-0.80762 -0.40104,-1.22132 -0.15625,-1.90625 0.25339,-0.70898 0.5725,-1.09805 0.9375,-0.96875 l 1.875,0.6875 c 0.0529,-0.21998 0.12303,-0.42855 0.21875,-0.625 l -1.875,-0.8125 c -0.40985,-0.17809 -0.50967,-0.48047 -0.15625,-1.1875 0.39027,-0.78065 0.66697,-1.07726 1.34375,-1.34375 0.70055,-0.27586 1.20087,-0.29739 1.34375,0.0625 l 0.75,1.90625 c 0.17927,-0.0814 0.36568,-0.14554 0.5625,-0.1875 l -0.59375,-2 c -0.13037,-0.42743 0.0139,-0.68527 0.78125,-0.875 0.42364,-0.10473 0.74466,-0.1426 1.03125,-0.125 z" style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#bebebe;fill:#000000;fill-opacity:1;stroke:none;stroke-width:5.61250019;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans" ns2:nodetypes="ssscscscsccsscccscccccsccccccccccccc"/>
        <ns0:path ns2:type="arc" style="color:#bebebe;fill:none;stroke:#000000;stroke-width:1.87825239;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path40342" ns2:cx="-30.94697" ns2:cy="239.58937" ns2:rx="2.8173785" ns2:ry="2.8173785" d="m -28.129591,239.58937 c 0,1.556 -1.261384,2.81738 -2.817379,2.81738 -1.555995,0 -2.817379,-1.26138 -2.817379,-2.81738 0,-1.55599 1.261384,-2.81738 2.817379,-2.81738 1.555995,0 2.817379,1.26139 2.817379,2.81738 z" transform="matrix(0.53240981,0,0,0.53240982,327.47647,95.44027)"/>
        <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:0.80000001;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible" d="m 318.96509,227.77445 c -0.0253,1.0815 -0.57608,2.26591 -2.37078,2.2245 -1.79469,-0.0413 -2.38091,-0.99117 -2.5307,-1.62378 C 313.91382,227.74255 313.69092,225 317.43304,223 c -1.43284,1.93104 1.56716,3.27382 1.53205,4.77445 z" id="path13227" ns2:nodetypes="szzcs"/>
      </ns0:g>
    </ns0:g>
    <ns0:g style="display:inline" id="g54146" ns1:label="haguichi" transform="matrix(2.680386,0,0,2.680386,-311.95426,-361.47556)">
      <ns0:rect transform="translate(241.0002,217)" y="18" x="-58" height="16" width="16" id="rect42965" style="fill:none;stroke:none"/>
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path54141" ns1:connector-curvature="0" d="m 193.569,236.00019 c -0.53334,0.0118 -1.06703,0.20368 -1.50255,0.58458 -1.40065,1.22494 -0.31275,2.49763 -1.53415,3.5658 -1.22144,1.0682 -2.30367,-0.20856 -3.70433,1.01639 l 0,0.002 c -0.31109,0.27206 -0.53556,0.60895 -0.67131,0.97299 -0.002,0.003 -0.002,0.005 -0.002,0.007 -0.0272,0.0741 -0.0508,0.14835 -0.0705,0.22438 -0.009,0.0337 -0.0188,0.0679 -0.0261,0.10182 -6.3e-4,0.005 -0.002,0.007 -0.002,0.0114 -0.0153,0.0719 -0.0266,0.14398 -0.0354,0.21683 -9e-5,4.9e-4 5e-5,0.002 0,0.002 -5.1e-4,0.005 -0.002,0.007 -0.002,0.0114 -0.005,0.0339 -0.007,0.0678 -0.0101,0.10182 -0.002,0.0257 -0.005,0.0516 -0.006,0.0774 -5.1e-4,0.0132 -0.002,0.0265 -0.002,0.0397 -1.2e-4,0.005 1e-4,0.008 0,0.0132 -6e-4,0.0343 -6e-4,0.0677 0,0.10182 2.5e-4,0.0174 0.002,0.0353 0.002,0.0527 0.002,0.0257 0.005,0.0516 0.006,0.0773 0.004,0.0379 0.007,0.0753 0.011,0.11313 8e-5,5e-4 -6e-5,0.002 0,0.002 0.009,0.0729 0.02,0.14499 0.0354,0.21687 6.1e-4,0.005 0.002,0.007 0.002,0.0114 0.007,0.0343 0.017,0.0679 0.0261,0.10182 0.0198,0.0761 0.0433,0.15036 0.0707,0.2244 0.002,0.003 0.002,0.005 0.002,0.007 0.13579,0.36407 0.36026,0.70094 0.67134,0.97302 l 0,0.002 c 1.40067,1.22494 2.48289,-0.0518 3.70431,1.01639 1.22142,1.06818 0.13352,2.34087 1.53417,3.56579 0.99548,0.87063 2.49799,0.75679 3.35656,-0.25265 0.85857,-1.00948 0.74817,-2.53305 -0.24735,-3.40366 -1.40063,-1.22495 -2.48287,0.0537 -3.70428,-1.01449 -0.61701,-0.53961 -0.64403,-1.13277 -0.70107,-1.74426 0.057,-0.61147 0.0842,-1.20464 0.70107,-1.74424 1.22141,-1.0682 2.30365,0.21044 3.70428,-1.0145 0.99552,-0.8706 1.10592,-2.39417 0.24735,-3.40364 -0.48294,-0.56782 -1.16828,-0.85234 -1.85402,-0.83724 z"/>
    </ns0:g>
    <ns0:g id="g30845" transform="matrix(0.67009649,0,0,0.67009649,131.52264,-246.54011)" ns1:label="file-roller">
      <ns0:path ns1:connector-curvature="0" ns1:original-d="m 346.83588,794.44498 -4.77297,15.55635 c 0,0 3.53553,10.78338 4.24264,10.25305 0.7071,-0.53033 24.39518,0 24.39518,0 l -0.88388,-14.31891 6.71751,-12.72792 z" ns1:path-effect="#path-effect30843" id="path30841" d="m 346.83588,794.44498 -4.77297,15.55635 c 0.18303,3.76817 1.70957,7.45731 4.24264,10.25305 3.07474,3.39357 7.61825,5.40802 12.19759,5.40802 4.57934,0 9.12285,-2.01445 12.19759,-5.40802 l -0.88388,-14.31891 6.71751,-12.72792 -29.69848,1.23743" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:g ns1:label="file-roller" id="g6474" style="display:inline" transform="matrix(3.9852721,0,0,3.9852721,-950.24365,71.174473)">
        <ns0:rect style="fill:none;stroke:none" id="rect6184" width="16" height="16" x="82" y="-42" transform="translate(241.0002,217)"/>
        <ns0:path ns1:connector-curvature="0" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:0.62873191;marker:none;visibility:visible;display:inline;overflow:visible" d="m 330.07659,187.00703 c 0,0 -2.91924,-0.0221 -3.10498,-0.0221 -0.18574,0 -0.26784,0.0324 -0.37159,-0.14741 -0.30689,-0.42982 -0.52143,-1.10364 -0.57752,-1.71708 -0.0109,-0.11882 -0.20696,-0.12631 -0.30151,-0.12683 L 323.15958,185 c -0.13341,0 -0.15695,0.24121 -0.15695,0.24121 -0.0519,1.89982 0.71945,4.7556 2.88858,4.74728 L 333.7812,190 c -2.67921,-0.16112 -2.63112,-1.34814 -2.84212,-2.47213 -0.18112,-0.35221 -0.25941,-0.52078 -0.5697,-0.52078 z" id="rect337" ns2:nodetypes="czcszccccccc" ns1:r_cx="true" ns1:r_cy="true"/>
        <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="path4320" d="m 332.0002,181.49621 2.5,0 c 3.80719,0 4.21897,8 0,8 l -2.9375,0" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.34051171;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 85.09375,-36 c -1.27743,0 -2.3125,2.02507 -2.3125,4.5 0,2.47494 1.03507,4.375 2.3125,4.375 0.0306,0 0.06355,-0.02925 0.09375,-0.03125 l 0,0.03125 8.812498,-0.875 c -1.8125,0 -3.062498,-1.098645 -3.062498,-3.5 0,-2.389424 1.03608,-3.5 3.062498,-3.5 l -1.585934,-0.996098 C 89.184425,-36.006039 85.09375,-36 85.09375,-36 z m 0.02344,0.992187 4.97656,0.0078 c 0.16968,2.66e-4 0.32247,0.18898 0.1875,0.375 -0.84239,1.515638 -0.897612,3.781759 -0.356694,5.569432 0,0.17445 -0.14283,0.3125 -0.3125,0.3125 l -5.048906,0.01386 c -0.16969,0 -0.25,-0.20055 -0.25,-0.375 -0.0858,-1.75606 -0.921312,-4.157719 0.585288,-5.841109 0,0 0.04901,-0.06277 0.218752,-0.0625 z" transform="translate(241.0002,217)" id="path5472" ns1:connector-curvature="0" ns2:nodetypes="csscccsccccsccccccsc"/>
        <ns0:path ns1:connector-curvature="0" style="fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none" d="m 330.00832,177 c -0.39473,0 -0.70961,0.17025 -0.88958,0.46259 l -2.28241,3.68924 -0.14046,0.27756 0.30433,0 1.10135,0 0.11704,0 0.0469,-0.10414 1.4538,-2.17057 c 0.0363,-0.0581 0.15888,-0.15034 0.28091,-0.15034 l 7.3961,0.003 c 0.0786,-0.005 0.079,0.10987 0.079,0.10987 l -2.87252,5.72088 -0.0937,0.16191 0.16385,0.0926 0.0698,0.70127 0.6942,0.36803 0.0936,-0.1619 3.46967,-7 c 0.13852,-0.23162 0.005,-1.3902 -0.10814,-1.59514 -0.12605,-0.22734 -0.3837,-0.41187 -0.71398,-0.40478 l -8.16989,0 z" id="path5477" ns2:nodetypes="cccccccccccccccccccsccc"/>
        <ns0:path transform="matrix(0.49627604,0,0,0.49230822,318.11937,169.76921)" ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path6840" ns2:cx="33.78125" ns2:cy="31.953125" ns2:rx="1.78125" ns2:ry="3.046875" d="M 35.5625,31.953125 C 35.5625,33.635868 34.765007,35 33.78125,35 32.797493,35 32,33.635868 32,31.953125 c 0,-1.682743 0.797493,-3.046875 1.78125,-3.046875 0.983757,0 1.78125,1.364132 1.78125,3.046875 z"/>
      </ns0:g>
    </ns0:g>
    <ns0:g transform="matrix(2.0102895,0,0,2.0102895,-304.991,-47.656345)" style="fill:#ffffff;fill-opacity:1;display:inline" id="g11071" ns1:label="seahorse">
      <ns0:path ns2:type="inkscape:offset" ns1:radius="0" ns1:original="M 247.40625 195.84375 C 245.19711 195.84375 243.40625 197.53552 243.40625 199.625 C 243.40625 201.16882 244.37959 202.50551 245.78125 203.09375 L 245.78125 203.84375 L 246.40625 203.84375 L 247.40625 204.84375 L 246.40625 205.84375 L 246.40625 206.84375 L 247.21875 207.84375 L 246.40625 208.3125 L 246.40625 208.75 L 247.40625 209.84375 L 248.40625 209.84375 L 249.40625 208.84375 L 249.40625 203.34375 C 249.25 203.28905 249.25295 203.3131 249.25 203.3125 C 247.98051 202.69626 247.0195 201.56142 246.625 200.1875 C 245.94432 200.1269 245.40625 199.53967 245.40625 198.84375 C 245.40625 198.15905 245.92881 197.607 246.59375 197.53125 C 246.76114 196.91261 247.02987 196.34211 247.40625 195.84375 z " ns4:href="#path11032" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3.33333325;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path30857" ns1:href="#path11032" d="m 247.40625,195.84375 c -2.20914,0 -4,1.69177 -4,3.78125 0,1.54382 0.97334,2.88051 2.375,3.46875 l 0,0.75 0.625,0 1,1 -1,1 0,1 0.8125,1 -0.8125,0.46875 0,0.4375 1,1.09375 1,0 1,-1 0,-5.5 c -0.15625,-0.0547 -0.1533,-0.0307 -0.15625,-0.0312 -1.26949,-0.61624 -2.2305,-1.75108 -2.625,-3.125 -0.68068,-0.0606 -1.21875,-0.64783 -1.21875,-1.34375 0,-0.6847 0.52256,-1.23675 1.1875,-1.3125 0.16739,-0.61864 0.43612,-1.18914 0.8125,-1.6875 z"/>
      <ns0:path ns2:type="inkscape:offset" ns1:radius="0" ns1:original="M 251.28125 195 C 250.18606 195 249.08641 195.40659 248.25 196.1875 C 247.4136 196.96841 247 197.97576 247 199 C 247 200.02424 247.4136 201.03159 248.25 201.8125 C 249.48924 202.96951 251.30794 203.24474 252.84375 202.6875 L 257.28125 207 L 258.5625 207 L 259 206.59375 L 259 204.75 L 258.25 204 L 257.5 204 L 256.75 202.5 L 256 202.5 L 256 201 L 255.25 200.4375 C 255.84684 199.0036 255.55173 197.34452 254.3125 196.1875 C 253.47609 195.40659 252.37644 195 251.28125 195 z M 250.5 196 C 251.32843 196 252 196.67157 252 197.5 C 252 198.32843 251.32843 199 250.5 199 C 249.67157 199 249 198.32843 249 197.5 C 249 196.67157 249.67157 196 250.5 196 z " ns4:href="#path234" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3.33333325;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path30855" ns1:href="#path234" d="m 251.28125,195 c -1.09519,0 -2.19484,0.40659 -3.03125,1.1875 -0.8364,0.78091 -1.25,1.78826 -1.25,2.8125 0,1.02424 0.4136,2.03159 1.25,2.8125 1.23924,1.15701 3.05794,1.43224 4.59375,0.875 l 4.4375,4.3125 1.28125,0 0.4375,-0.40625 0,-1.84375 -0.75,-0.75 -0.75,0 -0.75,-1.5 -0.75,0 0,-1.5 -0.75,-0.5625 c 0.59684,-1.4339 0.30173,-3.09298 -0.9375,-4.25 C 253.47609,195.40659 252.37644,195 251.28125,195 z M 250.5,196 c 0.82843,0 1.5,0.67157 1.5,1.5 0,0.82843 -0.67157,1.5 -1.5,1.5 -0.82843,0 -1.5,-0.67157 -1.5,-1.5 0,-0.82843 0.67157,-1.5 1.5,-1.5 z"/>
      <ns0:path ns1:connector-curvature="0" id="path234" d="m 251.28145,195 c -1.09519,0 -2.19484,0.40659 -3.03125,1.1875 -0.8364,0.78091 -1.25,1.78826 -1.25,2.8125 0,1.02424 0.4136,2.03159 1.25,2.8125 1.23924,1.15701 3.05794,1.43224 4.59375,0.875 l 4.4375,4.3125 1.28125,0 0.4375,-0.40625 0,-1.84375 -0.75,-0.75 -0.75,0 -0.75,-1.5 -0.75,0 0,-1.5 -0.75,-0.5625 c 0.59684,-1.4339 0.30173,-3.09298 -0.9375,-4.25 C 253.47629,195.40659 252.37664,195 251.28145,195 z m -0.78125,1 c 0.82843,0 1.5,0.67157 1.5,1.5 0,0.82843 -0.67157,1.5 -1.5,1.5 -0.82843,0 -1.5,-0.67157 -1.5,-1.5 0,-0.82843 0.67157,-1.5 1.5,-1.5 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="csccccccccccccccccscc" ns1:connector-curvature="0" id="path11032" d="m 247.41685,195.83334 c -2.20914,0 -4,1.69177 -4,3.78125 0,1.54382 0.97334,2.88051 2.375,3.46875 l 0,0.75 0.625,0 1,1 -1,1 0,1 0.81152,1 -0.81152,0.48614 0,0.4342 1,1.07966 1,0 1,-1 0,0 0,-5.47656 c -0.15625,-0.0547 -0.1533,-0.0541 -0.15625,-0.0547 -1.26949,-0.61624 -2.2305,-1.75108 -2.625,-3.125 -0.68068,-0.0606 -1.21875,-0.64783 -1.21875,-1.34375 0,-0.6847 0.52256,-1.23675 1.1875,-1.3125 0.16739,-0.61864 0.43612,-1.18914 0.8125,-1.6875 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:g>
    <ns0:g transform="matrix(0.67009649,0,0,0.67009649,112.52867,-18.739367)" id="g30934">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6.24000025;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path30936" ns2:cx="413" ns2:cy="560.86218" ns2:rx="29.5" ns2:ry="29.5" d="m 442.5,560.86218 c 0,16.2924 -13.2076,29.5 -29.5,29.5 -16.2924,0 -29.5,-13.2076 -29.5,-29.5 0,-16.2924 13.2076,-29.5 29.5,-29.5 16.2924,0 29.5,13.2076 29.5,29.5 z" transform="matrix(0.96153846,0,0,0.96153846,133.63462,24.821622)"/>
      <ns0:path ns2:nodetypes="sccccccccccsccccscccccscccccccccccccccccccccccccccs" ns1:connector-curvature="0" id="path159-6-3" d="m 538.58035,543.84408 c -1.47456,-0.0645 -2.22819,0.0972 -2.21708,0.11066 0.0213,0.0285 6.13645,1.15986 7.20553,2.66049 0,0 -2.55107,0.0248 -5.09929,0.77601 -0.11531,0.0356 9.36682,1.17492 11.30712,10.8637 0,0 -1.0413,-2.284 -2.32796,-2.66051 0.84613,2.62977 0.5841,7.71838 -0.22171,10.19858 -0.10357,0.3189 -0.18623,-1.37501 -1.77366,-2.10625 0.5084,3.72199 -0.0214,9.57 -2.54966,11.19628 -0.19685,0.12664 1.55879,-5.84933 0.33242,-3.54732 -7.32057,11.46674 -15.98026,4.65062 -19.51035,2.21709 2.8333,0.7093 6.38645,0.24971 7.5381,-0.55428 1.75846,-1.2279 2.83489,-2.09673 3.76902,-1.88453 0.93373,0.21321 1.50118,-0.81354 0.776,-1.66279 -0.726,-0.85097 -2.49267,-1.96774 -4.8776,-1.33028 -1.68195,0.45006 -3.69122,1.9251 -6.87295,0 -2.71442,-1.64308 -2.37942,-2.48105 -2.37942,-3.33116 0,-0.85057 0.75869,-2.09674 2.10624,-1.88455 0.30187,0.0475 0.53472,0.0318 0.66512,0 0.65565,0.1497 1.26793,0.34196 1.88454,0.66512 0.0285,-0.79494 -0.10361,-3.0984 -0.55427,-4.36363 0.0376,0.0141 0.1025,0.0389 0.11065,0 0.13622,-0.62741 3.74164,-0.65222 4.87362,-2.11573 0.72381,-0.93514 0.49922,-2.82663 0.49922,-2.82663 l -3.54732,0 c -1.85719,0.008 -3.44958,-2.66355 -3.59881,-3.03896 0.40594,-2.22052 1.72443,-2.97804 3.59881,-4.05571 -1.41,-0.0107 -0.66942,0 -3.54736,0 -1.87562,0 -3.00521,1.28266 -3.59878,1.94947 -2.48519,-0.58837 -4.90045,-0.89487 -6.5998,-0.21603 -0.78485,-0.81378 -1.40488,-2.8398 -1.49655,-5.28064 0,0 -4.27402,2.62017 -3.82444,9.04969 -0.008,0.52869 -0.17701,0.75728 -0.2217,1.10855 -0.46333,0.81039 -0.55091,1.43637 -0.44341,1.33023 -0.23273,0.4834 -0.54596,1.00753 -0.776,1.66282 -0.0528,0.12841 -0.17557,0.16424 -0.22169,0.33239 -0.0318,0.11422 0.008,0.22631 0,0.3324 -0.40838,1.28055 -0.76324,3.48503 -1.10855,5.47216 0,0 0.44073,-1.82421 1.10855,-3.14424 -0.55478,1.92808 -0.9298,5.49744 -0.66512,9.68465 0,0 0.0533,-0.72468 0.22169,-1.77366 0.16495,2.84146 0.91966,6.12753 2.99306,9.75515 5.1845,9.07231 13.80792,13.08558 22.83596,12.30482 1.57912,-0.10501 3.17978,-0.38432 4.76672,-0.77601 21.03296,-5.195 18.73433,-31.14975 18.73433,-31.14975 l -0.55426,3.8799 c 0,0 -0.85656,-7.09386 -1.88451,-9.75515 -1.57545,-4.07792 -2.21254,-4.10751 -2.21709,-4.1016 1.05511,2.73945 0.77598,4.21244 0.77598,4.21244 0,0 -1.81902,-5.10598 -6.76209,-6.7621 -2.92707,-0.98019 -5.17669,-1.37661 -6.65125,-1.44109 z" style="fill:#ffffff;fill-opacity:1;stroke:none;display:inline"/>
    </ns0:g>
    <ns0:g transform="matrix(0.67009649,0,0,0.67009649,152.16814,-192.18383)" id="g24776" ns1:label="documents">
      <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:7;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 608.17584,693.39936 -29.90154,9.20048 9.20047,28.43782 29.69243,-9.20047 z" id="path24774" ns1:connector-curvature="0"/>
      <ns0:rect y="687.36218" x="573" height="64" width="64" id="rect24747" style="color:#000000;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cccccc" ns1:connector-curvature="0" id="path21570" d="m 590.85066,695.9724 0,48.284 39.75057,0 0,-39.53456 -9.0735,-8.74944 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:5;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns1:connector-curvature="0" id="path24751" d="m 609.19489,730.79208 11.94524,-1.63633 -3.09102,-20.75399 m -12.80011,-8.22934 -19.02884,2.84563 4.39113,30.31973" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:nodetypes="cccccc"/>
      <ns0:path ns1:connector-curvature="0" id="path24749" d="m 608.17584,693.39936 -29.90154,9.20048 9.20047,28.43782 29.69243,-9.20047 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path style="color:#000000;fill:none;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 598.29097,704.40685 0,12.82105 -2.46912,2.89508 -2.82186,-3.30866 0,-26.05569 7.05464,0 0,4.5494" id="path24783" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:g id="g21476" transform="matrix(0.81617665,0,0,0.80644993,63.591961,-281.82582)">
      <ns0:path transform="translate(0,1)" d="m 587.53125,767.40625 c -0.26729,0.0807 -0.50363,0.24975 -0.6875,0.46875 -0.38334,0.45681 -0.3789,1.10005 -0.125,1.5625 l 0,0.0312 2.65625,4.75 c 0.006,0.0104 0.0677,0.14068 -0.21875,0.5625 -0.28416,0.41855 -0.82303,0.92507 -1.53125,1.3125 -0.71838,0.39296 -1.44476,0.57816 -1.9375,0.59375 -0.50359,0.0159 -0.61959,-0.084 -0.625,-0.0937 l -2.65625,-4.8125 c -0.23595,-0.42259 -0.5908,-0.66231 -1.0625,-0.71875 -0.47057,-0.0563 -0.917,0.0997 -1.21875,0.4375 -0.26765,0.28835 -0.29177,0.53808 -0.3125,0.625 -0.5566,2.43849 -0.31757,5.15779 0.8125,7.1875 1.47521,2.64964 4.46237,3.90403 7.40625,3.53125 0.94685,0.33714 2.28201,1.09453 3.90625,2.71875 l 21.78125,21.78125 c 1.39665,1.39664 2.14638,2.54682 2.5625,3.4375 -0.32625,1.59456 -0.18326,3.27342 0.65625,4.78125 1.12913,2.02805 3.31661,3.69814 5.6875,4.53125 0.5817,0.21597 1.2118,-0.057 1.53125,-0.4375 0.3358,-0.40018 0.44649,-1.03152 0.15625,-1.5625 l 0,-0.0312 -2.6875,-4.75 c -0.006,-0.0103 -0.0677,-0.14056 0.21875,-0.5625 0.28419,-0.41856 0.82305,-0.9251 1.53125,-1.3125 0.71836,-0.39296 1.44473,-0.57816 1.9375,-0.59375 0.50374,-0.0159 0.61963,0.0841 0.625,0.0937 l 2.6875,4.8125 c 0.18246,0.32683 0.54474,0.66054 1.03125,0.71875 0.4707,0.0563 0.91738,-0.10032 1.21875,-0.4375 0.14746,-0.15886 0.2689,-0.31116 0.34375,-0.625 0.55658,-2.43848 0.31758,-5.15778 -0.8125,-7.1875 -1.4849,-2.66704 -4.50588,-3.92395 -7.46875,-3.53125 -0.93069,-0.36018 -2.19003,-1.12753 -3.8125,-2.75 l -21.8125,-21.78125 c -1.42497,-1.42496 -2.14052,-2.60945 -2.53125,-3.53125 0.29383,-1.55756 0.13256,-3.18333 -0.6875,-4.65625 -1.12914,-2.02804 -3.31661,-3.69814 -5.6875,-4.53125 -0.30664,-0.11383 -0.60771,-0.11199 -0.875,-0.0312 z" id="path21474" style="fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none;display:inline;enable-background:new" ns1:original="M 588.09375 768.3125 C 587.90788 768.2435 587.68848 768.3187 587.5625 768.46875 C 587.43654 768.61885 587.43186 768.82821 587.53125 769 L 590.1875 773.78125 C 590.42649 774.21053 590.28855 774.74951 589.90625 775.3125 C 589.5204 775.88084 588.88577 776.45589 588.0625 776.90625 C 587.23906 777.35668 586.40789 777.6032 585.71875 777.625 C 585.03368 777.6467 584.48962 777.46164 584.25 777.03125 L 581.59375 772.21875 C 581.51915 772.08514 581.37003 771.98685 581.21875 771.96875 C 581.06756 771.95067 580.91313 772.01234 580.8125 772.125 C 580.7582 772.1835 580.73736 772.26573 580.71875 772.34375 C 580.21076 774.56927 580.45978 777.11893 581.4375 778.875 C 582.77274 781.27324 585.53961 782.4144 588.25 781.9375 C 589.3589 782.3154 590.84761 783.16013 592.59375 784.90625 L 614.375 806.6875 C 615.90831 808.2208 616.76356 809.52893 617.21875 810.5625 C 616.80593 812.07436 616.94915 813.68661 617.75 815.125 C 618.72729 816.88032 620.77161 818.45767 622.9375 819.21875 C 623.12335 819.28775 623.31154 819.21255 623.4375 819.0625 C 623.56346 818.91239 623.5995 818.70304 623.5 818.53125 L 620.8125 813.75 C 620.5735 813.32072 620.71157 812.78175 621.09375 812.21875 C 621.47961 811.65044 622.11423 811.07535 622.9375 810.625 C 623.76093 810.17457 624.5921 809.92806 625.28125 809.90625 C 625.96631 809.88465 626.51038 810.0696 626.75 810.5 L 629.4375 815.3125 C 629.5121 815.44613 629.62997 815.5444 629.78125 815.5625 C 629.93254 815.5806 630.08685 815.51886 630.1875 815.40625 C 630.2418 815.34775 630.29389 815.26553 630.3125 815.1875 C 630.82047 812.96198 630.57147 810.41232 629.59375 808.65625 C 628.25228 806.24683 625.44116 805.09933 622.71875 805.59375 C 621.62933 805.18921 620.20481 804.32981 618.46875 802.59375 L 596.65625 780.8125 C 595.08217 779.23843 594.26835 777.87647 593.84375 776.8125 C 594.20648 775.34392 594.05519 773.79633 593.28125 772.40625 C 592.30395 770.65093 590.25964 769.07357 588.09375 768.3125 z " ns1:radius="0.92327356" ns2:type="inkscape:offset"/>
      <ns0:path d="m 623.15625,772.84375 a 3.1822988,3.1822988 0 0 0 -1.625,0.59375 l -2.75,1.9375 a 3.1822988,3.1822988 0 0 0 -0.71875,0.71875 l -1.75,2.375 -16,16.03125 a 3.1822988,3.1822988 0 0 0 -0.0312,0 3.1822988,3.1822988 0 0 0 -3.9375,1.21875 c 0,0 -0.63972,1.00096 -1.375,2.09375 -0.36764,0.54639 -0.77526,1.09883 -1.09375,1.53125 -0.31849,0.43242 -0.72144,0.83829 -0.40625,0.5625 0.24157,-0.21138 -1.15819,0.79124 -2.40625,1.59375 -1.24806,0.80251 -2.54175,1.59011 -3.65625,2.625 -1.15536,1.07283 -2.36395,2.62613 -3.5625,4.125 -1.19855,1.49887 -2.21875,2.8125 -2.21875,2.8125 a 3.1822988,3.1822988 0 0 0 -0.5625,2.71875 c 0,0 0.14195,0.52076 0.375,1.15625 0.23305,0.63549 0.48875,1.41396 1.3125,2.375 1.24969,1.45797 2.18219,1.52412 2.96875,1.78125 0.78656,0.25713 1.46875,0.40625 1.46875,0.40625 a 3.1822988,3.1822988 0 0 0 2.59375,-0.625 c 0,0 1.47716,-1.16436 3.125,-2.53125 1.64784,-1.36689 3.3037,-2.69177 4.4375,-4 1.02245,-1.17975 1.72819,-2.48113 2.40625,-3.625 0.67806,-1.14387 1.47783,-2.20996 1.28125,-2.03125 0.1192,-0.10836 1.15946,-0.815 2,-1.3125 0.84054,-0.4975 1.5625,-0.875 1.5625,-0.875 a 3.1822988,3.1822988 0 0 0 1.375,-4.15625 l -0.0625,-0.0937 15.96875,-16 2.375,-1.625 a 3.1822988,3.1822988 0 0 0 0.78125,-0.71875 l 2.125,-2.875 A 3.1822988,3.1822988 0 0 0 626.71875,774.75 L 625.5,773.65625 a 3.1822988,3.1822988 0 0 0 -2.34375,-0.8125 z" id="path21472" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:4;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:original="M 623.375 776.03125 L 620.625 777.96875 L 618.6875 780.59375 L 600.84375 798.4375 L 599.03125 797.40625 C 599.03125 797.40625 596.37755 801.59934 595.5625 802.3125 C 594.74746 803.02567 590.98883 805.1443 589.5625 806.46875 C 588.13617 807.7932 584.15625 813 584.15625 813 C 584.15625 813 584.54497 814.53684 585.15625 815.25 C 585.76754 815.96317 587.8125 816.375 587.8125 816.375 C 587.8125 816.375 593.61305 811.77821 594.9375 810.25 C 596.26195 808.72179 597.78557 805.36256 598.90625 804.34375 C 600.02694 803.32495 603.09375 801.6875 603.09375 801.6875 L 602.09375 799.5625 L 619.8125 781.8125 L 622.46875 780 L 624.59375 777.125 L 623.375 776.03125 z " ns1:radius="3.1819806" ns2:type="inkscape:offset"/>
    </ns0:g>
    <ns0:g transform="matrix(0.67009649,0,0,0.67009649,174.50084,-225.78817)" id="g25797">
      <ns0:rect y="530.34058" x="673.07727" height="64" width="64" id="rect25795" style="color:#000000;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:rect ry="2.4805617" rx="2.4805617" y="539.61224" x="717.70361" height="15.50351" width="10.852457" id="rect25714" style="color:#000000;fill:#edf3fb;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:rect ry="2.4805617" rx="2.4805617" y="552.41345" x="718.67584" height="15.193439" width="11.782667" id="rect25716" style="color:#000000;fill:#edf3fb;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:rect ry="2.277133" rx="2.488415" y="565.36646" x="716.48029" height="16.793856" width="15.863646" id="rect25718" style="color:#000000;fill:#edf3fb;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-linecap:square;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:rect ry="2.4960177" rx="2.4805617" y="534.2077" x="678.05804" height="57.096397" width="48.060883" id="rect25712" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:4;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path style="font-size:23.55376053px;font-style:normal;font-weight:normal;fill:url(#radialGradient25776);fill-opacity:1;stroke:none;display:inline;enable-background:new;font-family:Bitstream Vera Sans" id="path5099" d="m 700.43477,563.41392 c -2e-5,1.41414 0.28918,2.52934 0.86758,3.34562 0.5895,0.81629 1.38479,1.22443 2.38587,1.22443 0.98992,0 1.77964,-0.40814 2.36918,-1.22443 0.58949,-0.82777 0.88425,-1.94298 0.88427,-3.34562 -2e-5,-1.39112 -0.30034,-2.48908 -0.90096,-3.29388 -0.58953,-0.81627 -1.38482,-1.22442 -2.38586,-1.22443 -0.97883,10e-6 -1.763,0.40816 -2.3525,1.22443 -0.5784,0.8048 -0.8676,1.90276 -0.86758,3.29388 m 6.84059,5.19088 c -0.33371,0.81629 -0.87317,1.45437 -1.61839,1.91425 -0.73413,0.44838 -1.59615,0.67258 -2.58607,0.67258 -1.91316,0 -3.47037,-0.71282 -4.67162,-2.13844 -1.19017,-1.43712 -1.78524,-3.30538 -1.78523,-5.60478 -10e-6,-2.29938 0.60062,-4.16764 1.80191,-5.60477 1.20126,-1.43711 2.7529,-2.15567 4.65494,-2.15569 0.98992,2e-5 1.85194,0.22996 2.58607,0.68982 0.74522,0.4599 1.28468,1.09798 1.61839,1.91425 l 0,-2.25916 3.48703,0 0,11.95111 c 1.37922,-0.21844 2.4637,-0.90251 3.25345,-2.05221 0.7897,-1.16119 1.18456,-2.6443 1.18459,-4.44933 -3e-5,-1.14969 -0.16131,-2.22465 -0.48385,-3.2249 -0.32259,-1.01172 -0.81199,-1.93723 -1.46822,-2.77652 -1.0567,-1.40262 -2.38033,-2.48333 -3.97088,-3.24215 -1.57947,-0.75878 -3.2924,-1.13818 -5.13878,-1.1382 -1.29028,2e-5 -2.52492,0.17823 -3.70393,0.53461 -1.17904,0.34493 -2.26909,0.85655 -3.27014,1.53485 -1.6462,1.12672 -2.93089,2.58683 -3.85408,4.38034 -0.91209,1.78205 -1.36813,3.71354 -1.36812,5.79448 -10e-6,1.71306 0.29475,3.32263 0.88427,4.82873 0.60063,1.49461 1.46265,2.81676 2.58608,3.96645 1.11228,1.12671 2.38585,1.98323 3.82071,2.56958 1.44597,0.59784 2.98649,0.89676 4.62157,0.89676 1.40147,0 2.80296,-0.27018 4.20446,-0.81053 1.40147,-0.54036 2.59718,-1.27042 3.58714,-2.19018 l 1.78523,2.79377 c -1.39039,1.1152 -2.90867,1.96598 -4.55484,2.55233 -1.63508,0.59783 -3.29796,0.89675 -4.98862,0.89676 -2.05775,-10e-6 -3.9987,-0.37941 -5.82284,-1.1382 -1.82417,-0.74731 -3.44811,-1.83952 -4.87184,-3.27664 -1.42373,-1.43712 -2.50822,-3.09843 -3.25345,-4.98394 -0.74523,-1.89699 -1.11785,-3.93196 -1.11785,-6.10489 0,-2.09244 0.37818,-4.08716 1.13454,-5.98418 0.75635,-1.89698 1.83527,-3.56404 3.23676,-5.00118 1.40148,-1.42561 3.03098,-2.52931 4.88852,-3.31113 1.86864,-0.78177 3.80402,-1.17266 5.80616,-1.17269 2.49151,3e-5 4.75502,0.49439 6.79053,1.48311 2.03547,0.97726 3.73728,2.39139 5.10542,4.24238 0.83419,1.12673 1.46264,2.35115 1.88534,3.67328 0.43376,1.31067 0.65066,2.69031 0.65069,4.13892 -3e-5,3.11569 -0.90655,5.5358 -2.71955,7.26034 -1.81307,1.72454 -4.37133,2.58682 -7.67481,2.58682 l -0.65069,0 0,-2.65581" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:g transform="matrix(0.67009649,0,0,0.67009649,174.50084,-209.98391)" id="g4666">
      <ns0:rect style="color:#000000;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25795-7" width="64" height="64" x="673.07727" y="610.34058"/>
      <ns0:path ns1:connector-curvature="0" id="path11079-0-4" d="m 681.5,619.875 c -0.57222,0 -1,0.32189 -1,1.03125 l 0,12 -0.65625,0 c -0.78383,0 -1.3115,0.72566 -1.3125,1.21875 l 0,5.96875 c -0.0287,9.14657 -0.23851,24.78125 2.0625,24.78125 l 48.78125,0 c 2.15452,0 2.129,-10.76297 2.125,-23.78125 l 0,-12 c -2e-4,-0.73962 -0.52865,-1.21875 -1.3125,-1.21875 l -0.6875,0 0,-1.78125 c 0,-0.78365 -0.47994,-1.1875 -1.09375,-1.1875 l -23.03125,0 c -0.41474,0 -1.06817,-0.0817 -1.59375,-0.6875 l -3.21875,-3.6875 c -0.44856,-0.51696 -1.01194,-0.65625 -1.46875,-0.65625 l -17.59375,0 z" style="fill:#ffffff;stroke:#000000;stroke-width:6;stroke-miterlimit:4;stroke-dasharray:none;display:inline;enable-background:new"/>
      <ns0:path ns1:connector-curvature="0" style="fill:#ffffff;stroke:#000000;stroke-width:0.99999994;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 680.74059,634.34791 11.84823,-0.005 c 0.94491,-3.4e-4 1.6868,-0.44095 2.14934,-1.03839 l 1.7296,-2.54936 c 0.35778,-0.52736 0.98464,-0.89347 1.7096,-0.89347 l 29.11052,0 c 0.72469,0 1.20761,0.43981 1.20779,1.09948 l 0.004,10.71456 c 0.004,11.61098 0.0282,21.18618 -1.96361,21.18618 l -45.09853,0 c -2.12734,0 -1.94893,-13.92337 -1.92236,-22.08119 l 0.0183,-5.33415 c 9.2e-4,-0.43979 0.48313,-1.09949 1.20779,-1.09949 l -2e-5,0 0,0 z" id="path9590-3-9" ns2:nodetypes="czzszczzcczzcccc" ns1:r_cx="true" ns1:r_cy="true"/>
      <ns0:path ns2:nodetypes="ccccccccscccccscccccccccccccccccccccccccccccc" ns1:connector-curvature="0" id="path4642-7" d="m 695.55752,654.98582 0,0.0311 c -0.4677,1.49346 0.005,3.02317 1.2735,3.9459 1.26886,0.92308 2.88563,0.90628 4.16216,0 l 0.0311,0 m 3.97579,-2.85845 3.9758,2.85845 0.0311,0 c 1.27653,0.90628 2.8933,0.92308 4.16216,0 1.26837,-0.92273 1.7412,-2.45244 1.2735,-3.9459 l 0,-0.0311 -1.45986,-4.62944 3.94473,-2.95166 c 0.0105,-0.0103 0.0208,-0.0206 0.0311,-0.0311 1.24619,-0.94625 1.70614,-2.46118 1.21138,-3.94589 -0.4914,-1.47462 -1.7733,-2.40193 -3.32352,-2.42347 l -0.0311,0 -4.8455,-0.0621 -1.58411,-4.66051 c -0.52351,-1.55658 -1.9412,-2.44576 -3.572,-2.36132 -0.0135,7e-4 -0.0175,-0.0319 -0.0311,-0.0311 -0.0109,6.8e-4 -0.0202,-7.7e-4 -0.0311,0 l 0,0.0311 c -1.46379,0.0996 -2.66507,0.96378 -3.13715,2.36132 l -1.58411,4.66051 -4.8455,0.0621 -0.0311,0 c -1.55022,0.0215 -2.83212,0.94885 -3.32352,2.42347 m 1.21138,3.94589 c 0.0102,0.0105 0.0206,0.0208 0.0311,0.0311 l 3.94473,2.95166 m -0.52803,-5.37518 5.03186,-0.0621 c 0.81384,-0.009 1.59337,-0.56808 1.86366,-1.33601 l 1.61516,-4.78479 1.61517,4.78479 c 0.27029,0.76793 1.04982,1.32675 1.86366,1.33601 l 5.03186,0.0621 -4.03791,2.98273 c -0.66144,0.49192 -0.96185,1.41954 -0.71441,2.20597 l 1.52199,4.81586 -4.1311,-2.92059 m -3.94271,1.16241 -2.4869,1.75818 0.85496,-2.70524" style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans"/>
    </ns0:g>
    <ns0:g transform="matrix(0.67009649,0,0,0.67009649,174.52673,-194.17964)" id="g6123">
      <ns0:rect y="690.34058" x="673.07727" height="64" width="64" id="rect25795-7-5" style="color:#000000;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path transform="matrix(0.40741882,0,0,0.40741883,664.18837,680.72101)" d="m 156.62415,104.66175 c 0,35.24482 -28.57157,63.81639 -63.816388,63.81639 -35.244817,0 -63.816387,-28.57157 -63.816387,-63.81639 0,-35.244817 28.57157,-63.816386 63.816387,-63.816386 35.244818,0 63.816388,28.571569 63.816388,63.816386 z" ns2:ry="63.816387" ns2:rx="63.816387" ns2:cy="104.66175" ns2:cx="92.807762" id="path6667-6-2-12" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:14.72686195;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      <ns0:path ns1:connector-curvature="0" id="path7720-2-1" d="m 710.46875,704.78125 -1.9375,0.375 c 0.0625,0.11195 0.13497,0.22584 0.1875,0.34375 0.0624,0.15499 0.0983,0.30982 0.125,0.46875 l 1.75,-0.34375 c 0.002,-0.2907 -0.0388,-0.56504 -0.125,-0.84375 z m -0.59375,2.6875 -5.6875,1.125 c 0.0164,0.0716 0.0152,0.14801 0.0625,0.21875 0.20906,0.26525 0.4914,0.45539 0.8125,0.5625 0.3989,0.1117 0.80813,0.1306 1.21875,0.0625 0.32194,-0.0616 0.61943,-0.17094 0.90625,-0.28125 0.0983,0.16409 0.18646,0.31731 0.25,0.5 l 1.78125,-0.34375 c -0.01,-0.18199 -0.0404,-0.35253 -0.0937,-0.53125 -0.0633,-0.17844 -0.12791,-0.36734 -0.21875,-0.53125 0.0931,-0.061 0.18594,-0.12384 0.28125,-0.1875 0.25529,-0.16838 0.48247,-0.37063 0.6875,-0.59375 z m -17.625,1.8125 c -0.21805,0.0211 -0.43995,0.0253 -0.65625,0.0625 -0.28877,0.0521 -0.56881,0.12024 -0.84375,0.21875 l 1.5,-0.28125 z m 5.59375,0.5625 -3.65625,0.71875 c 0.40941,0.0527 0.81295,0.11112 1.21875,0.1875 0.57027,0.10995 1.1316,0.23638 1.6875,0.40625 0.34704,0.10747 0.69027,0.21904 1.03125,0.34375 L 701,710.9375 c -0.24067,-0.10682 -0.47513,-0.21225 -0.71875,-0.3125 -0.51659,-0.20561 -1.06395,-0.39407 -1.59375,-0.5625 -0.27013,-0.085 -0.53761,-0.15189 -0.8125,-0.21875 l -0.0312,0 z m 10.78125,1.3125 -1.4375,0.28125 c -0.0863,0.14499 -0.19861,0.27686 -0.3125,0.40625 -0.23848,0.0631 -0.4735,0.12204 -0.71875,0.15625 -0.48804,0.0599 -0.98011,0.0372 -1.46875,0 -0.0721,-0.006 -0.14697,-0.0229 -0.21875,-0.0312 l -3.4375,0.6875 c 0.17993,0.0566 0.37943,0.11012 0.5625,0.15625 0.50519,0.13229 1.0106,0.26 1.53125,0.3125 0.49613,0.0435 0.9712,0.0771 1.46875,0.0312 0.47317,-0.0539 0.9647,-0.12418 1.40625,-0.3125 0.93196,-0.43611 1.90532,-0.93512 2.625,-1.6875 z m -20.53125,0.625 -1.28125,0.25 c -0.24068,0.22959 -0.46806,0.46903 -0.6875,0.71875 -0.35421,0.40137 -0.68602,0.85894 -0.96875,1.3125 -0.005,0.008 0.005,0.023 0,0.0312 l 1.5,-0.3125 c 0.0892,-0.17113 0.17644,-0.33711 0.28125,-0.5 0.28843,-0.44411 0.57904,-0.89015 0.9375,-1.28125 0.0677,-0.0735 0.14966,-0.14653 0.21875,-0.21875 z m -2.1875,3.875 -1.5625,0.3125 c -0.13233,0.41903 -0.24496,0.81519 -0.3125,1.25 -0.078,0.4566 -0.0746,0.92222 0,1.375 l 1.84375,-0.375 c -0.0367,-0.12153 -0.0724,-0.24784 -0.0937,-0.375 -0.0853,-0.48665 -0.12265,-0.97965 -0.0312,-1.46875 0.0424,-0.24379 0.0944,-0.47968 0.15625,-0.71875 z m 20.53125,2.03125 c -0.25316,-0.007 -0.49782,0.0133 -0.75,0.0625 -0.57941,0.12425 -1.16369,0.32392 -1.71875,0.53125 -0.5515,0.19686 -1.10559,0.36326 -1.65625,0.5625 -0.5704,0.20525 -1.14724,0.39165 -1.71875,0.59375 -0.58489,0.20429 -1.16859,0.41094 -1.75,0.625 -0.58843,0.1984 -1.15521,0.41474 -1.75,0.59375 -0.5678,0.17938 -1.14139,0.35354 -1.71875,0.5 -0.57936,0.14378 -1.15903,0.25825 -1.75,0.34375 -0.59117,0.0799 -1.18485,0.13575 -1.78125,0.0937 -0.5739,-0.0418 -1.16097,-0.10507 -1.71875,-0.25 -0.53155,-0.14128 -1.05749,-0.31096 -1.5625,-0.53125 -0.45958,-0.20396 -0.9312,-0.4286 -1.34375,-0.71875 -0.14392,-0.10887 -0.27474,-0.22171 -0.40625,-0.34375 l -2.125,0.4375 c 0.25151,0.36048 0.5603,0.66714 0.90625,0.9375 0.41726,0.30747 0.90518,0.53584 1.375,0.75 0.51017,0.22917 1.02436,0.38256 1.5625,0.53125 0.33269,0.0921 0.69014,0.16947 1.03125,0.21875 l 8.875,-1.78125 c 0.21747,-0.0767 0.43867,-0.14234 0.65625,-0.21875 0.57261,-0.1987 1.14675,-0.39327 1.71875,-0.59375 0.55057,-0.19933 1.10347,-0.40071 1.65625,-0.59375 0.55272,-0.20407 1.11459,-0.36195 1.6875,-0.5 0.48459,-0.1143 0.98025,-0.10995 1.46875,-0.0312 0.3162,0.0595 0.58242,0.20191 0.84375,0.375 l 2.25,-0.46875 c -0.10291,-0.13819 -0.21204,-0.25799 -0.34375,-0.375 -0.34889,-0.2952 -0.73744,-0.54892 -1.1875,-0.65625 -0.25008,-0.0518 -0.49684,-0.087 -0.75,-0.0937 z m 2.71875,2.75 -1.6875,0.34375 c 0.0143,0.2075 -0.006,0.41853 -0.0625,0.625 -0.12437,0.3718 -0.35134,0.66641 -0.59375,0.96875 -0.20282,0.23322 -0.44569,0.43256 -0.6875,0.625 -0.4527,0.17856 -0.93281,0.32776 -1.40625,0.4375 -0.54877,0.12303 -1.09898,0.20855 -1.65625,0.28125 -0.58832,0.0746 -1.1588,0.11145 -1.75,0.15625 -0.61418,0.0353 -1.23125,0.0996 -1.84375,0.15625 -0.63083,0.0599 -1.28131,0.14686 -1.90625,0.25 -0.61928,0.0946 -1.20582,0.21971 -1.8125,0.375 -0.56225,0.14178 -1.12619,0.32913 -1.65625,0.5625 -1.02661,0.51137 -2.0914,1.02536 -2.90625,1.84375 -0.32296,0.33483 -0.55582,0.72359 -0.71875,1.15625 -0.1334,0.36827 -0.15305,0.7727 -0.0937,1.15625 0.076,0.37396 0.30798,0.66269 0.5625,0.9375 0.2797,0.30185 0.61449,0.54547 0.96875,0.75 0.41117,0.22785 0.83205,0.36811 1.28125,0.5 0.50675,0.14314 1.04306,0.23 1.5625,0.3125 0.53389,0.0705 1.06934,0.15874 1.59375,0.28125 0.46747,0.11375 0.90188,0.31347 1.3125,0.5625 0.35307,0.22548 0.62703,0.52059 0.84375,0.875 0.17247,0.29981 0.241,0.62849 0.25,0.96875 -0.008,0.34225 -0.13365,0.67123 -0.21875,1 -0.11248,0.38597 -0.1646,0.7872 -0.1875,1.1875 -0.0146,0.42495 0.0615,0.83792 0.15625,1.25 0.10047,0.41223 0.2997,0.804 0.53125,1.15625 0.2495,0.37418 0.57806,0.67313 0.9375,0.9375 0.37996,0.25377 0.765,0.49962 1.125,0.78125 0.18012,0.13603 0.34354,0.27578 0.5,0.4375 l 1.625,-1 c -0.16043,-0.1703 -0.31344,-0.32623 -0.5,-0.46875 -0.36101,-0.28434 -0.73856,-0.56365 -1.125,-0.8125 -0.34589,-0.24478 -0.66849,-0.5197 -0.90625,-0.875 -0.22024,-0.33231 -0.4099,-0.67129 -0.5,-1.0625 -0.0875,-0.39606 -0.15,-0.8114 -0.125,-1.21875 0.0304,-0.39015 0.10986,-0.77989 0.21875,-1.15625 0.0884,-0.34452 0.16715,-0.67208 0.15625,-1.03125 -0.0218,-0.3704 -0.0932,-0.73727 -0.28125,-1.0625 -0.23174,-0.37896 -0.5036,-0.71868 -0.875,-0.96875 -0.41985,-0.26897 -0.89136,-0.46771 -1.375,-0.59375 -0.52622,-0.13199 -1.05547,-0.21315 -1.59375,-0.28125 -0.51396,-0.0778 -1.02859,-0.17792 -1.53125,-0.3125 -0.43872,-0.12211 -0.87663,-0.25594 -1.28125,-0.46875 -0.34253,-0.18835 -0.66829,-0.40036 -0.9375,-0.6875 -0.23289,-0.24177 -0.41165,-0.50505 -0.46875,-0.84375 -0.0415,-0.35764 -0.0149,-0.7275 0.125,-1.0625 0.17905,-0.40887 0.42352,-0.75408 0.75,-1.0625 0.0637,-0.0581 0.11556,-0.0883 0.15625,-0.125 0.3537,-0.14423 0.72214,-0.28009 1.09375,-0.375 0.60163,-0.16499 1.19597,-0.30985 1.8125,-0.40625 0.62241,-0.1042 1.24689,-0.21705 1.875,-0.28125 0.61167,-0.0569 1.2301,-0.0933 1.84375,-0.125 0.5929,-0.0427 1.19092,-0.1169 1.78125,-0.1875 0.56027,-0.069 1.10344,-0.13409 1.65625,-0.25 0.51088,-0.11062 1.04195,-0.21951 1.53125,-0.40625 1.03351,-0.40842 1.99861,-0.98604 2.90625,-1.625 0.35165,-0.2749 0.6946,-0.5823 0.96875,-0.9375 0.24234,-0.32591 0.4652,-0.66147 0.5625,-1.0625 0.008,-0.0406 -0.006,-0.0844 0,-0.125 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:path style="color:#000000;fill:#000000;stroke:#000000;stroke-width:1;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 724.69874,693.95992 -12.90842,21.14191 c -0.62566,0.95205 1.17028,3.25354 4.01136,5.14051 2.8411,1.88696 5.65145,2.64484 6.27711,1.69279 L 736.359,701.70432 c 0.70908,-1.079 -1.32516,-3.68916 -4.54505,-5.82771 -3.21987,-2.13856 -6.40613,-2.99569 -7.11521,-1.91669 z" id="use6644-3-5-1" ns1:connector-curvature="0" ns2:nodetypes="ccsccsc"/>
      <ns0:path clip-path="none" ns2:nodetypes="csccscc" ns1:connector-curvature="0" id="path10325-06" d="m -898.25,55.250002 c -15.56651,-1.966347 -62.00971,11.685352 -77,3.75 -25.102,-13.288176 -40.5049,-17.66697 -68.5,-22.5 l 0.25,-3.25 c 0,0 32.5143,-6.411419 49.65541,-13.160732 9.73303,-3.832377 70.48998,0.745769 93.93124,1.87132 5.24,8.346471 5.9344,22.192941 1.66335,33.289412 z" style="fill:#ffffff;stroke:#000000;stroke-width:4.84004307;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline;enable-background:new" transform="matrix(0.11388834,-0.17238628,0.17238628,0.11388834,814.27804,556.97443)"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path10341-6" d="m 708.74248,728.98369 -7.17426,11.81686" style="fill:#000000;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline;enable-background:new"/>
      <ns0:path transform="matrix(0.07775427,-0.1176922,0.19503281,0.12884995,753.69289,648.34237)" d="m -644.52783,30.592316 c 0,0.97631 -2.29523,1.767767 -5.12653,1.767767 -2.8313,0 -5.12652,-0.791457 -5.12652,-1.767767 0,-0.976311 2.29522,-1.767767 5.12652,-1.767767 2.8313,0 5.12653,0.791456 5.12653,1.767767 z" ns2:ry="1.767767" ns2:rx="5.126524" ns2:cy="30.592316" ns2:cx="-649.65436" id="path10343-0" style="color:#000000;fill:url(#radialGradient10861-2);fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:8.26067448;stroke-miterlimit:4;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
    </ns0:g>
    <ns0:g transform="matrix(0.67009649,0,0,0.67009649,174.50084,-178.37538)" id="g6861">
      <ns0:rect style="color:#000000;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25795-7-5-8" width="64" height="64" x="673.07727" y="770.34058"/>
      <ns0:path ns2:nodetypes="sscccccccsssccscccccsss" ns1:connector-curvature="0" id="path6383" d="m 686.28125,787.34375 c -0.65368,0 -1.18343,0.13167 -1.71875,0.375 -0.53532,0.24333 -1.14286,0.55598 -1.6875,1.5 l -5.40625,12.375 c -0.20139,0.34906 -0.49281,0.94134 -0.5,1.90625 l -0.0312,0 0,0.0937 0,9.375 c -5e-5,0.0104 -5e-5,0.0208 0,0.0312 0.007,0.88499 0.45524,1.95206 1.21875,2.59375 0.76351,0.64169 1.64947,0.84375 2.34375,0.84375 l 24.75,0 c 0.74787,0 1.52633,-0.28532 2.1875,-0.75 0.012,-0.008 0.0193,-0.0226 0.0312,-0.0312 0.95903,-0.52423 1.59375,-1.59454 1.59375,-2.6875 l 0,-9.46875 c 0.004,-0.30606 -0.0384,-0.61268 -0.125,-0.90625 -0.003,-0.0188 0.004,-0.0439 0,-0.0625 l -1.8125,-12.34375 c -0.002,-0.0106 0.002,-0.0207 0,-0.0312 -0.24038,-1.19295 -1.01232,-1.93766 -1.65625,-2.3125 -0.64961,-0.37814 -1.2838,-0.5 -1.9375,-0.5 z" style="color:#000000;fill:#ffffff;stroke:#000000;stroke-width:6;stroke-linejoin:round;stroke-miterlimit:4;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path6453-7" d="m 681,804.86218 6.125,0" style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path6453-7-3" d="m 681,808.86218 2.625,0" style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1"/>
      <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="path6453-7-3-2" d="m 681,810.86218 3.75,0 m 13.125,0 4.125,0" style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1"/>
      <ns0:path ns2:nodetypes="ccccc" ns1:connector-curvature="0" id="path6578" d="m 686.34375,791.46875 -4.875,11.84375 22.34375,0 -1.625,-11.84375 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.62994266;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path6453-7-3-27" d="m 701.375,806.86218 4.625,0" style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1"/>
      <ns0:path ns2:nodetypes="sssssssss" ns1:connector-curvature="0" id="path6828" d="m 699.71875,778.375 c -2.01271,0 -3.6875,1.68933 -3.6875,3.6875 l 0,36.59375 c 0,1.99817 1.67479,3.6875 3.6875,3.6875 l 25.5625,0 c 2.01271,0 3.6875,-1.68933 3.6875,-3.6875 l 0,-36.59375 c 0,-1.99817 -1.67479,-3.6875 -3.6875,-3.6875 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6;stroke-miterlimit:4;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(4,0)"/>
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 706.74999,790.36218 c -0.41421,0 -0.75,0.27996 -0.75,0.62532 0,0.73067 1.21875,0.92723 1.5,1.77173 0.28125,-0.8445 1.5,-1.04106 1.5,-1.77173 0,-0.34536 -0.33579,-0.62532 -0.75,-0.62532 -0.41421,0 -0.75,0.27996 -0.75,0.62532 0,-0.34536 -0.33579,-0.62532 -0.75,-0.62532 z" id="path3904-7-8-4" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 714.24999,795.41805 c -1.24263,0 -2.25,0.99243 -2.25,2.21666 0,2.59012 3.65626,3.28691 4.50001,6.28053 0.84374,-2.99362 4.5,-3.69041 4.5,-6.28053 0,-1.22423 -1.00737,-2.21666 -2.25,-2.21666 -1.24265,0 -2.25,0.99243 -2.25,2.21666 0,-1.22423 -1.00736,-2.21666 -2.25001,-2.21666 z" id="path3904-1-9-2" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 726.25,810.36218 c 0.41421,0 0.75,-0.27996 0.75,-0.62532 0,-0.73067 -1.21875,-0.92723 -1.5,-1.77173 -0.28125,0.8445 -1.5,1.04106 -1.5,1.77173 0,0.34536 0.33579,0.62532 0.75,0.62532 0.41421,0 0.75,-0.27996 0.75,-0.62532 0,0.34536 0.33579,0.62532 0.75,0.62532 z" id="path3904-7-8-6-5" ns1:connector-curvature="0"/>
      <ns0:path style="opacity:0.7;color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 707.5,785.36218 c -0.831,0 -1.5,0.669 -1.5,1.5 l 0,0.5 0,1 0,1 1,0 0,-1 1,0 0,1 1,0 0,-1 0,-1 0,-0.5 c 0,-0.831 -0.669,-1.5 -1.5,-1.5 z m 0,1 c 0.277,0 0.5,0.223 0.5,0.5 l 0,0.5 -1,0 0,-0.5 c 0,-0.277 0.223,-0.5 0.5,-0.5 z" id="rect6648-9" ns1:connector-curvature="0"/>
      <ns0:path style="opacity:0.7;color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 725.5,815.36218 c -0.831,0 -1.5,-0.669 -1.5,-1.5 l 0,-0.5 0,-1 0,-1 1,0 0,1 1,0 0,-1 1,0 0,1 0,1 0,0.5 c 0,0.831 -0.669,1.5 -1.5,1.5 z m 0,-1 c 0.277,0 0.5,-0.223 0.5,-0.5 l 0,-0.5 -1,0 0,0.5 c 0,0.277 0.223,0.5 0.5,0.5 z" id="rect6648-1-7" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:g id="g7498" mask="url(#mask8354)" transform="translate(58,176)">
      <ns0:g id="g5606" transform="matrix(0.67009649,0,0,0.67009649,67.09785,-193.37936)">
        <ns0:rect y="840.34058" x="583.07727" height="64" width="64" id="rect25795-7-5-8-7-4" style="color:#000000;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
        <ns0:path style="fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6;stroke-miterlimit:4;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 596.96875,846.34375 c -4.91834,0 -9,4.08165 -9,9 l 0,24.0625 c 0,4.91835 4.08166,9 9,9 l 18.1875,0 -0.0215,10.19988 13.61527,-10.19988 4.28125,0 c 4.91835,0 9,-4.08165 9,-9 l 0,-24.0625 c 0,-4.91835 -4.08165,-9 -9,-9 z" id="path5513" ns1:connector-curvature="0" ns2:nodetypes="sssscccsssss"/>
        <ns0:path ns1:connector-curvature="0" id="rect3165-6-2-1-6-6-5-0-0-2-2-5-2" d="m 621.2306,856.33486 -6.07584,5.97267 -5.8695,-5.97267 -9.13362,-0.0496 10.53844,10.48685 -10.84794,10.59003 8.82411,-0.10113 6.48851,-6.02427 6.12741,6.02427 8.87569,-0.002 -10.53844,-10.48686 10.48686,-10.43527 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:nodetypes="ccccccccccccc"/>
      </ns0:g>
      <ns0:g id="g6852" transform="matrix(0.67009649,0,0,0.67009649,74.09785,-193.37936)">
        <ns0:g id="g6522" transform="matrix(1.2027105,0,0,1.2027105,-142.37053,-173.36379)">
          <ns0:path ns2:nodetypes="cccccccssssccssccccccc" ns1:connector-curvature="0" id="path3073-4" d="m 727,845.36218 -20.65625,0.125 0,29.78125 -3.03125,0.15625 -13.5,0 c -7.27846,1.78742 -8.44185,12.76551 -8.3125,17.875 l 1.21875,0 0,-0.125 c 0,-0.36674 0.29271,-1.15625 0.625,-1.15625 l 2.0625,0 c 0.33229,0 0.59375,0.78951 0.59375,1.15625 l 0,0.0937 16.625,0.125 c 0.0157,-0.35099 0.30293,-1 0.625,-1 l 1.8125,0 c 0.31275,0 0.62729,0.63222 0.65625,0.96875 l 0.75,0 c -0.17844,-2.58741 1.0253,-6.09883 1.6875,-8.53125 l 15.78125,-0.0625 -0.002,0 c 1.42089,0 3.00157,-2.23306 3.00157,-6.1875 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:#000000;stroke-width:4.98873138;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
          <ns0:path ns1:connector-curvature="0" ns2:nodetypes="ccsccscc" id="path4008-0" d="m 725.37635,847.0251 -17.46512,0.12614 0.0184,28.75142 c 0.002,3.18513 -1.04094,3.94707 -1.66979,4.53598 l 16.26018,4.18533 c 1.25753,0 2.80654,-2.19565 2.80654,-6.0516 l 0.0499,-31.54727 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible"/>
          <ns0:path ns1:connector-curvature="0" ns2:nodetypes="ccccc" id="path3230-9" d="m 690.2652,877.57803 25.35473,-0.38547 c 5.57574,0 3.68849,6.91996 9.38007,8.02751 0,0 -28.33503,-0.0651 -28.33503,-0.0651 l -6.39977,-7.57695 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible"/>
          <ns0:path ns2:type="inkscape:offset" ns1:radius="-0.61472619" ns1:original="M 134.375 28.46875 L 110.15625 28.5 C 103.12278 30.227252 102.125 40.8125 101.875 45.875 L 102.75 45.875 L 102.75 45.5625 C 102.75 45.208103 103.02264 44.9375 103.34375 44.9375 L 104.09375 44.9375 C 104.41486 44.9375 104.6875 45.208103 104.6875 45.5625 L 104.6875 45.84375 L 122.9375 45.65625 L 122.9375 45.5 C 122.9375 45.145603 123.21014 44.875 123.53125 44.875 L 124.28125 44.875 C 124.60236 44.875 124.875 45.145603 124.875 45.5 L 124.875 45.625 L 125.9375 45.625 C 125.9375 45.625 126.3763 30.848731 134.375 28.46875 z " ns4:href="#path3119" style="color:#000000;fill:#ffffff;stroke:url(#linearGradient6529);stroke-width:0.56242812;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:0.5624281, 2.24971244;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path3145-4" d="M 131.8125,29.09375 110.25,29.125 c -3.1975,0.819607 -5.06865,3.628614 -6.1875,7 -0.96869,2.918941 -1.27418,6.044683 -1.4375,8.5 0.2061,-0.169389 0.4359,-0.3125 0.71875,-0.3125 l 0.75,0 c 0.53432,0 0.90334,0.415856 1.0625,0.90625 L 122.5,45.03125 c 0.18962,-0.429042 0.54145,-0.78125 1.03125,-0.78125 l 0.75,0 c 0.47543,0 0.80282,0.340593 1,0.75 l 0.0937,0 c 0.0363,-0.775432 0.19634,-3.653053 1.1875,-7.21875 0.89893,-3.233921 2.48383,-6.727577 5.25,-8.6875 z" transform="matrix(1.0348322,0,0,1.0348322,575.76665,846.16023)" ns1:href="#path3119"/>
          <ns0:path style="fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 692.65558,875.19275 0.80847,0 c 0.34172,0 0.45532,0.0681 0.2587,0.1617 l -0.38806,0.19403 c -0.19662,0.0936 -0.62843,0.16169 -0.97015,0.16169 l -0.8408,0 c -0.34173,0 -0.45533,-0.0681 -0.25871,-0.16169 l 0.4204,-0.19403 c 0.19662,-0.0936 0.62843,-0.1617 0.97015,-0.1617 z m 15.49219,1.09951 0.80846,0 c 0.34172,0 0.48766,0.14071 0.29105,0.29105 l -0.42041,0.29105 c -0.19661,0.15034 -0.62843,0.2587 -0.97015,0.2587 l -0.80846,0 c -0.34173,0 -0.45533,-0.10836 -0.25871,-0.2587 l 0.38806,-0.29105 c 0.19662,-0.15034 0.62843,-0.29105 0.97016,-0.29105 z m -17.72354,0.0647 0.80846,0 c 0.34172,0 0.48766,0.1407 0.29105,0.29105 l -0.42041,0.29104 c -0.19661,0.15035 -0.62843,0.25871 -0.97015,0.25871 l -0.80846,0 c -0.34173,0 -0.45533,-0.10836 -0.25871,-0.25871 l 0.38806,-0.29104 c 0.19662,-0.15035 0.62843,-0.29105 0.97016,-0.29105 z m -2.00499,1.8433 0.80846,0 c 0.34172,0 0.45533,0.16478 0.25871,0.38806 l -0.4204,0.45274 c -0.19662,0.22327 -0.62843,0.4204 -0.97016,0.4204 l -0.80846,0 c -0.34172,0 -0.45533,-0.19713 -0.25871,-0.4204 l 0.38806,-0.45274 c 0.19662,-0.22328 0.66078,-0.38806 1.0025,-0.38806 z m 18.1116,0 0.80846,0 c 0.34173,0 0.45533,0.16478 0.25871,0.38806 l -0.4204,0.45274 c -0.19662,0.22328 -0.62843,0.4204 -0.97015,0.4204 l -0.80847,0 c -0.34172,0 -0.45532,-0.19712 -0.25871,-0.4204 l 0.38807,-0.45274 c 0.19662,-0.22328 0.66077,-0.38806 1.00249,-0.38806 z m -19.63151,2.06966 0.74378,0 c 0.34408,0 0.5001,0.22938 0.35573,0.48508 l -0.32339,0.58209 c -0.14437,0.25569 -0.5614,0.45274 -0.90548,0.45274 l -0.71144,0 c -0.34407,0 -0.5001,-0.19705 -0.35573,-0.45274 l 0.32339,-0.58209 c 0.14437,-0.2557 0.52907,-0.48508 0.87314,-0.48508 z m 17.98225,0.0647 0.8408,0 c 0.34407,0 0.50009,0.22938 0.35572,0.48507 l -0.29105,0.51742 c -0.14436,0.25569 -0.5614,0.45274 -0.90547,0.45274 l -0.80847,0 c -0.34407,0 -0.50009,-0.19705 -0.35572,-0.45274 l 0.29105,-0.51742 c 0.14437,-0.25569 0.52907,-0.48507 0.87314,-0.48507 z m -19.08176,2.36071 0.77612,0 c 0.32482,0 0.46728,0.25793 0.35573,0.58209 l -0.22637,0.67911 c -0.11156,0.32416 -0.45131,0.58209 -0.77613,0.58209 l -0.77612,0 c -0.32481,0 -0.49962,-0.25793 -0.38806,-0.58209 l 0.22637,-0.67911 c 0.11155,-0.32416 0.48365,-0.58209 0.80846,-0.58209 z m 17.91757,0 0.97016,0 c 0.32481,0 0.46727,0.25793 0.35572,0.58209 l -0.22637,0.67911 c -0.11156,0.32416 -0.45131,0.58209 -0.77612,0.58209 l -0.97016,0 c -0.32481,0 -0.49962,-0.25793 -0.38806,-0.58209 l 0.22637,-0.67911 c 0.11155,-0.32416 0.48365,-0.58209 0.80846,-0.58209 z m -18.82305,2.97514 0.8408,0 c 0.35131,0 0.59386,0.27407 0.51742,0.61443 l -0.16169,0.67911 c -0.0765,0.34037 -0.42482,0.61443 -0.77613,0.61443 l -0.8408,0 c -0.3513,0 -0.56152,-0.27406 -0.48508,-0.61443 l 0.1617,-0.67911 c 0.0765,-0.34036 0.39248,-0.61443 0.74378,-0.61443 z m 18.1116,0 0.8408,0 c 0.35131,0 0.59386,0.27407 0.51742,0.61443 l -0.16169,0.67911 c -0.0765,0.34037 -0.42482,0.61443 -0.77613,0.61443 l -0.8408,0 c -0.3513,0 -0.56152,-0.27406 -0.48507,-0.61443 l 0.16169,-0.67911 c 0.0765,-0.34036 0.39248,-0.61443 0.74378,-0.61443 z m -18.532,2.9428 0.80846,0 c 0.3323,0 0.5821,0.31237 0.5821,0.67911 l 0,0.74379 c 0,0.36674 -0.2498,0.64677 -0.5821,0.64677 l -0.80846,0 c -0.33229,0 -0.61443,-0.28003 -0.61443,-0.64677 l 0,-0.74379 c 0,-0.36674 0.28214,-0.67911 0.61443,-0.67911 z m 18.1116,0 0.80847,0 c 0.33229,0 0.58209,0.31237 0.58209,0.67911 l 0,0.74379 c 0,0.36674 -0.2498,0.64677 -0.58209,0.64677 l -0.80847,0 c -0.33229,0 -0.61443,-0.28003 -0.61443,-0.64677 l 0,-0.74379 c 0,-0.36674 0.28214,-0.67911 0.61443,-0.67911 z" id="path7433" ns1:connector-curvature="0" ns2:nodetypes="ssccssccsssccssccsssccssccsssccssccsssccssccsssccssccsssccssccsssccssccsssccssccsssccssccsssccssccsssssssssssssssssss"/>
        </ns0:g>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531" width="2.0123537" height="2" x="710" y="846.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0" width="2.0123537" height="2" x="710" y="850.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0-5" width="2.0123537" height="2" x="710" y="854.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-9" width="2.0123537" height="2" x="710" y="858.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0-2" width="2.0123537" height="2" x="710" y="862.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0-5-4" width="2.0123537" height="2" x="710" y="866.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-9-1" width="2.0123537" height="2" x="710" y="870.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0-2-0" width="2.0123537" height="2" x="710" y="874.36218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-6" width="2.0123537" height="2" x="726.99384" y="846.61218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0-6" width="2.0123537" height="2" x="726.99384" y="850.61218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0-5-8" width="2.0123537" height="2" x="726.99384" y="854.61218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-9-12" width="2.0123537" height="2" x="726.99384" y="858.61218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.69999999;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6531-0-2-2" width="2.0123537" height="2" x="726.99384" y="862.61218" rx="0.35355338" ry="0.35355338"/>
        <ns0:rect style="color:#000000;fill:none;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25795-7-5-8-7-4-3" width="64" height="64" x="673.07727" y="840.34058"/>
      </ns0:g>
      <ns0:g id="g7363" transform="matrix(0.66014572,0,0,0.66014572,-96.53681,20.72842)">
        <ns0:path transform="matrix(0.96153846,0,0,0.96153846,133.63462,24.821622)" d="m 442.5,560.86218 c 0,16.2924 -13.2076,29.5 -29.5,29.5 -16.2924,0 -29.5,-13.2076 -29.5,-29.5 0,-16.2924 13.2076,-29.5 29.5,-29.5 16.2924,0 29.5,13.2076 29.5,29.5 z" ns2:ry="29.5" ns2:rx="29.5" ns2:cy="560.86218" ns2:cx="413" id="path7365" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:6.24000025;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
        <ns0:g ns1:transform-center-y="34.344176" ns1:transform-center-x="10.791579" transform="matrix(0.31132618,-0.02705993,0.02705993,0.31132618,416.64896,523.26137)" id="g7367" style="display:inline;enable-background:new">
          <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 353.89029,162.43914 c -0.8148,0 -1.50438,0.49404 -1.81876,1.1916 -0.01,0.0203 -0.0127,0.0426 -0.0207,0.0626 l -29.75544,65.2389 0.0208,0.0206 c -0.10568,0.19141 -0.16726,0.41393 -0.16726,0.64802 0,0.73893 0.59899,1.33796 1.33791,1.33796 0.51126,0 0.94549,-0.28936 1.17075,-0.71078 l 0.0626,-0.10453 c 0.0143,-0.0341 0.0303,-0.0692 0.0421,-0.10453 l 30.75888,-64.40268 0.0421,-0.0421 c 0.0962,-0.14236 0.15163,-0.31565 0.20906,-0.48082 0.007,-0.0144 0.0159,-0.0275 0.0207,-0.0421 0.0622,-0.19398 0.10452,-0.39144 0.10452,-0.60625 0,-1.10833 -0.89849,-2.00688 -2.00693,-2.00688 z" id="path7369" ns1:connector-curvature="0" ns2:nodetypes="cccccsscccccccscc"/>
        </ns0:g>
        <ns0:g transform="matrix(0.3118804,0.01966854,-0.01966854,0.3118804,489.29329,510.78749)" ns1:transform-center-y="-21.161415" ns1:transform-center-x="-4.9738117" id="g7371" style="display:inline;enable-background:new">
          <ns0:g style="fill:#000000;fill-opacity:1;stroke:none" id="g7373" clip-path="url(#clipPath6996-2)" transform="translate(-110,0)">
            <ns0:path ns2:nodetypes="csccccccccscccccc" ns1:connector-curvature="0" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 290.13291,107.02249 c -0.52316,-1.95241 -2.52999,-3.11107 -4.4824,-2.58791 -0.96349,0.25817 -1.73966,0.87495 -2.20981,1.67092 l -0.0311,-0.0182 -33.7284,55.3598 c -0.10281,0.17003 -0.19825,0.34177 -0.28097,0.52259 l 0.008,0.0245 -0.28755,0.49803 0.0621,0.0359 c -0.28822,0.89781 -0.33736,1.8833 -0.0752,2.86186 0.72658,2.71169 3.51384,4.32089 6.22554,3.5943 1.43104,-0.38344 2.54552,-1.34541 3.18122,-2.56271 l 0.0311,0.0182 0.28402,-0.7076 31.0997,-56.23417 c 0.34119,-0.74663 0.43404,-1.62082 0.20495,-2.47567 z" id="path7375"/>
            <ns0:path id="path7377" d="m 290.13291,107.02249 c -0.52316,-1.95241 -2.52999,-3.11107 -4.4824,-2.58791 -0.96349,0.25817 -1.73966,0.87495 -2.20981,1.67092 l -0.0311,-0.0182 -33.7284,55.3598 c -0.10281,0.17003 -0.19825,0.34177 -0.28097,0.52259 l 0.008,0.0245 -0.28755,0.49803 0.0621,0.0359 c -0.28822,0.89781 -0.33736,1.8833 -0.0752,2.86186 0.72658,2.71169 3.51384,4.32089 6.22554,3.5943 1.43104,-0.38344 2.54552,-1.34541 3.18122,-2.56271 l 0.0311,0.0182 0.28402,-0.7076 31.0997,-56.23417 c 0.34119,-0.74663 0.43404,-1.62082 0.20495,-2.47567 z" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0" ns2:nodetypes="csccccccccscccccc"/>
          </ns0:g>
          <ns0:g id="g7379" clip-path="url(#clipPath7139-5)" transform="translate(-140,0)">
            <ns0:path ns1:connector-curvature="0" id="path7381" d="m 257,136.25 c -2.48528,0 -4.5,2.01472 -4.5,4.5 0,1.22647 0.48552,2.34456 1.28125,3.15625 l -0.0312,0.0312 25.75,24.375 c 0.16907,0.17638 0.34266,0.34436 0.53125,0.5 l 0.0312,0 0.5,0.5 0.0625,-0.0625 c 0.97462,0.62799 2.12939,1 3.375,1 3.45178,0 6.25,-2.79822 6.25,-6.25 0,-1.82164 -0.78781,-3.45138 -2.03125,-4.59375 l 0.0312,-0.0312 -0.75,-0.5625 -27.625,-21.53125 C 259.09687,136.63839 258.08816,136.25 257,136.25 z" style="color:#000000;fill:url(#linearGradient7395);fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
            <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 257,136.25 c -2.48528,0 -4.5,2.01472 -4.5,4.5 0,1.22647 0.48552,2.34456 1.28125,3.15625 l -0.0312,0.0312 25.75,24.375 c 0.16907,0.17638 0.34266,0.34436 0.53125,0.5 l 0.0312,0 0.5,0.5 0.0625,-0.0625 c 0.97462,0.62799 2.12939,1 3.375,1 3.45178,0 6.25,-2.79822 6.25,-6.25 0,-1.82164 -0.78781,-3.45138 -2.03125,-4.59375 l 0.0312,-0.0312 -0.75,-0.5625 -27.625,-21.53125 C 259.09687,136.63839 258.08816,136.25 257,136.25 z" id="path7383" ns1:connector-curvature="0"/>
          </ns0:g>
          <ns0:path transform="matrix(0.26022189,0,0,0.26022189,-0.6833974,-113.79205)" d="m 600,1068 c 0,24.3005 -19.69947,44 -44,44 -24.30053,0 -44,-19.6995 -44,-44 0,-24.3005 19.69947,-44 44,-44 24.30053,0 44,19.6995 44,44 z" ns2:ry="44" ns2:rx="44" ns2:cy="1068" ns2:cx="556" id="path7385" style="fill:#000000;fill-opacity:1;stroke:none;display:inline;enable-background:new" ns2:type="arc"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g7387" transform="matrix(0.66014572,0,0,0.66014572,8.2967858,19.19907)">
        <ns0:path ns1:connector-curvature="0" ns1:original-d="m 478.18096,537.76522 -18.73833,18.73833 14.84924,8.30851 18.03123,-5.83363 0,-6.36397 z" ns1:path-effect="#path-effect30869" id="path7389" d="m 478.18096,537.76522 -18.73833,18.73833 14.84924,8.30851 18.03123,-5.83363 0,-6.36397 -14.14214,-14.84924" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:10;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:g transform="matrix(3.7500031,0,0,3.7521005,-830.66729,-1500.7311)" ns1:label="inkscape" id="g7391" style="display:inline">
          <ns0:path ns1:connector-curvature="0" id="path7393" d="m 348.94707,543.0052 c -0.45398,0 -0.8959,0.16964 -1.24379,0.52861 l -6.18785,6.37443 c -0.34097,0.35183 -0.52184,0.81575 -0.52861,1.27489 -1e-4,0.007 0,0.0234 0,0.031 -6e-5,1.36608 3.65031,0.04 3.98012,1.71022 0.17851,0.90395 -1.99006,0.48981 -1.99006,1.39927 0,1.06688 3.06954,0.3332 3.94903,1.21269 0.36128,0.87948 -1.17511,0.73753 -0.90174,1.55474 0.5152,0.53164 1.67415,0.23016 1.89678,1.08832 0.25429,0.98026 1.91986,0.81115 2.89181,0.0931 0.5152,-0.53162 -0.79505,-0.77436 -0.27984,-1.30597 0.51519,-0.53163 3.05996,-0.4241 3.07838,-1.58584 -0.24319,-0.72981 -1.19805,-0.84765 -1.21272,-1.71021 -0.0512,-0.73049 0.78195,-0.51683 3.42043,-1.2438 1.05503,-0.49441 1.09237,-0.75739 1.08832,-1.2127 -8e-5,-0.009 0,-0.0214 0,-0.031 -0.006,-0.45914 -0.21875,-0.92306 -0.5597,-1.27489 l -6.15676,-6.37443 c -0.34788,-0.35901 -0.78981,-0.52861 -1.2438,-0.52861 z m 0.12437,1.33708 c 0.46755,0.004 1.74874,1.58409 2.89182,2.76743 0.32152,0.42998 -0.12437,0.87065 -0.12437,0.87065 l -2.3943,-1.30598 -1.05723,1.43037 -0.93282,-1.39928 -0.55972,2.17664 -1.64802,-0.99504 0.43533,-0.55969 2.58086,-2.64306 c 0.19795,-0.2011 0.34952,-0.3456 0.80845,-0.34204 z m 7.08961,9.57719 c -0.12574,-0.004 -0.25257,0.006 -0.34204,0.031 -0.16865,0.0486 -0.96755,0.077 -0.90174,0.68409 0.72383,0.3034 1.82743,0.54491 1.95897,-0.0621 0.0988,-0.4552 -0.3379,-0.63905 -0.71519,-0.65297 z m -12.34461,2.02114 c -0.0702,0.008 -0.11793,0.036 -0.18656,0.0621 -0.54894,0.20872 -0.91708,0.64774 -0.40424,0.83956 0.51291,0.1918 0.85636,-0.0109 1.30597,-0.24876 0.44967,-0.23797 0.43675,-0.28133 0.40424,-0.37313 -0.0623,0.0125 -0.47121,-0.24203 -0.90174,-0.27987 -0.0717,-0.006 -0.14746,-0.008 -0.21767,0 z" style="fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none"/>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g7397" transform="matrix(0.67009649,0,0,0.67009649,-111.80834,-39.09348)">
        <ns0:path d="m 415.5,624.875 c -3.80438,0 -6.875,0.82143 -6.875,1.84375 l 0,36.1875 c 0,1.02233 3.07062,1.84375 6.875,1.84375 l 39.4375,0 c 3.80437,0 6.875,-0.82142 6.875,-1.84375 l 0,-36.1875 c 0,-1.02232 -3.07063,-1.84375 -6.875,-1.84375 l -7.375,0 -0.0937,0.46875 -9.25,0.0312 -0.125,-0.5 -22.59375,0 z" ns1:href="#rect19224" id="path7399" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:12;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns4:href="#rect19224" ns1:original="M 415.5 624.875 C 411.69562 624.875 408.625 625.69643 408.625 626.71875 L 408.625 662.90625 C 408.625 663.92858 411.69562 664.75 415.5 664.75 L 454.9375 664.75 C 458.74187 664.75 461.8125 663.92858 461.8125 662.90625 L 461.8125 626.71875 C 461.8125 625.69643 458.74187 624.875 454.9375 624.875 L 447.5625 624.875 L 447.46875 625.34375 L 438.21875 625.375 L 438.09375 624.875 L 415.5 624.875 z " ns1:radius="0" ns2:type="inkscape:offset"/>
        <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:6;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 415.50021,624.86773 22.58279,0.008 0.13613,0.48403 9.24186,-0.0303 0.10588,-0.46134 7.38138,0 c 3.80437,0 6.8671,0.82302 6.8671,1.84534 l 0,36.18087 c 0,1.02233 -3.06273,1.84535 -6.8671,1.84535 l -39.44804,0 c -3.80438,0 -6.86711,-0.82302 -6.86711,-1.84535 l 0,-36.18087 c 0,-1.02232 3.06273,-1.84534 6.86711,-1.84534 z" id="path7401" ns1:connector-curvature="0" ns2:nodetypes="sccccssssssss"/>
        <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:4.13201761;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter52127);enable-background:new" d="m 112.3125,52.53125 c -9.91951,0 -17.96875,2.850005 -17.96875,6.34375 0,1.933127 2.464014,3.652134 6.34375,4.8125 L 98.375,66.5 106,68 l 2.875,-2.53125 c 0.6345,0.02389 1.53499,0.21875 2.1875,0.21875 11.16951,0 19.1875,-3.318755 19.1875,-6.8125 0,-3.493745 -8.01799,-6.34375 -17.9375,-6.34375 z" transform="matrix(0.24201252,0,0,0.24201252,397.84496,613.66803)" id="path7403" ns1:connector-curvature="0" ns2:nodetypes="ssccccsss"/>
        <ns0:g transform="matrix(0.37915538,0,0,0.37915538,374.62159,591.25572)" id="g7405">
          <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.55063653;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter16757-8);enable-background:new" d="m 153.25,84.866387 42,0 1.6875,9.258613 -43.75,0 z" id="path7407" ns1:connector-curvature="0" ns2:nodetypes="ccccc"/>
          <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.39318216;marker:none;visibility:visible;display:inline;overflow:visible;filter:url(#filter16757-8);enable-background:new" id="path7409" ns2:cx="182.6875" ns2:cy="87.5625" ns2:rx="3.4375" ns2:ry="1.5625" d="m 186.125,87.5625 c 0,0.862945 -1.53902,1.5625 -3.4375,1.5625 -1.89848,0 -3.4375,-0.699555 -3.4375,-1.5625 0,-0.862945 1.53902,-1.5625 3.4375,-1.5625 1.89848,0 3.4375,0.699555 3.4375,1.5625 z" transform="matrix(1.1740571,0,0,1.6705259,-40.505155,-57.027801)"/>
          <ns0:g clip-path="none" id="g7411" transform="matrix(-1,0,0.19314882,1,337.86402,0)">
            <ns0:path transform="matrix(1,0,0,0.92018529,0.25,7.5447954)" ns2:nodetypes="cscccsccc" ns1:connector-curvature="0" id="path7413" d="m 161.44607,93.616606 c 0,0 -0.78005,-0.459575 -0.73974,-0.90054 0.0572,-0.62659 -0.1991,-1.501402 1.21733,-1.474766 l 5.94382,-0.0055 -0.0833,-12.140633 -4.68188,-0.09685 c -3.45297,-0.07143 -3.18065,2.428014 -3.18065,2.428014 l -0.0623,12.190276 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.55063653;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" clip-path="none"/>
          </ns0:g>
          <ns0:g transform="translate(-6.10467,0)" id="g7415" clip-path="none">
            <ns0:path clip-path="none" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.55063653;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 161.44607,93.616606 c 0,0 -0.78005,-0.459575 -0.73974,-0.90054 0.0572,-0.62659 -0.1991,-1.501402 1.21733,-1.474766 l 5.94382,-0.0055 -0.0833,-12.140633 -4.68188,-0.09685 c -3.45297,-0.07143 -3.18065,2.428014 -3.18065,2.428014 l -0.0623,12.190276 z" id="path7417" ns1:connector-curvature="0" ns2:nodetypes="cscccsccc" transform="matrix(1,0,0,0.92018529,0,7.5447954)"/>
          </ns0:g>
        </ns0:g>
        <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:4.01754808;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path7419" ns2:cx="69.125" ns2:cy="83.5" ns2:rx="18.625" ns2:ry="6.5" d="M 87.75,83.5 C 87.75,87.089851 79.411303,90 69.125,90 58.838697,90 50.5,87.089851 50.5,83.5 50.5,79.910149 58.838697,77 69.125,77 79.411303,77 87.75,79.910149 87.75,83.5 z" transform="matrix(0.2742272,0,0,0.22592655,436.28476,607.87482)"/>
        <ns0:g transform="matrix(0.26269733,0,0,0.26269733,398.17699,601.56142)" id="g7421">
          <ns0:path transform="matrix(0.73543852,0,0,0.73543852,47.808877,47.521858)" d="m 199.25,179.625 c 0,11.80509 -9.56991,21.375 -21.375,21.375 -11.80509,0 -21.375,-9.56991 -21.375,-21.375 0,-11.80509 9.56991,-21.375 21.375,-21.375 11.80509,0 21.375,9.56991 21.375,21.375 z" ns2:ry="21.375" ns2:rx="21.375" ns2:cy="179.625" ns2:cx="177.875" id="path7423" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.23782039;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
          <ns0:g id="g7425" transform="matrix(0.70175439,0,0,0.70175439,53.274123,53.572369)"/>
          <ns0:g id="g7427" clip-path="url(#clipPath15654)" transform="matrix(1.2642868,0,0,1.2642868,-370.38728,-93.77475)">
            <ns0:g id="g7429" transform="translate(0,6)"/>
            <ns0:g id="g7431" transform="translate(0,-3)">
              <ns0:path transform="matrix(0.82352941,0,0,1,76.213235,4)" d="m 446.75,218.9375 c 0,4.86701 -5.23267,8.8125 -11.6875,8.8125 -6.45483,0 -11.6875,-3.94549 -11.6875,-8.8125 0,-4.86701 5.23267,-8.8125 11.6875,-8.8125 6.45483,0 11.6875,3.94549 11.6875,8.8125 z" ns2:ry="8.8125" ns2:rx="11.6875" ns2:cy="218.9375" ns2:cx="435.0625" id="path7434" style="color:#000000;fill:#191025;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
              <ns0:path transform="matrix(0.66251783,0,0,0.88269156,146.26334,26.183217)" d="m 446.75,218.9375 c 0,4.86701 -5.23267,8.8125 -11.6875,8.8125 -6.45483,0 -11.6875,-3.94549 -11.6875,-8.8125 0,-4.86701 5.23267,-8.8125 11.6875,-8.8125 6.45483,0 11.6875,3.94549 11.6875,8.8125 z" ns2:ry="8.8125" ns2:rx="11.6875" ns2:cy="218.9375" ns2:cx="435.0625" id="path7436" style="color:#000000;fill:url(#radialGradient7468);fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
              <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path7438" ns2:cx="434.5" ns2:cy="218.5" ns2:rx="5.5" ns2:ry="5.5" d="m 440,218.5 c 0,3.03757 -2.46243,5.5 -5.5,5.5 -3.03757,0 -5.5,-2.46243 -5.5,-5.5 0,-3.03757 2.46243,-5.5 5.5,-5.5 3.03757,0 5.5,2.46243 5.5,5.5 z" transform="matrix(1.1363636,0,0,1.1363636,-59.25,-31.545455)"/>
              <ns0:path id="path7440" d="m 424.58196,217.89188 c -0.007,-0.13515 -0.0168,-0.26536 -0.0168,-0.40215 0,-4.53716 4.34257,-8.77776 9.62229,-8.77776 5.27973,0 9.4973,4.2406 9.4973,8.77776 0,0.13679 -0.009,0.267 -0.0168,0.40215 -0.2474,-4.34766 -4.48503,-6.62561 -9.60557,-6.62561 -5.12056,0 -9.23319,2.27795 -9.48059,6.62561 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns1:connector-curvature="0" ns2:nodetypes="cssscscc"/>
              <ns0:g id="g7442" transform="matrix(0.8813906,0,0,0.8813906,53.848934,25.653047)">
                <ns0:path transform="matrix(1.1582075,-0.27647923,0,1.1582075,-91.614292,75.799371)" d="m 452.75,224.25 c 0,1.51878 -1.45507,2.75 -3.25,2.75 -1.79493,0 -3.25,-1.23122 -3.25,-2.75 0,-1.51878 1.45507,-2.75 3.25,-2.75 1.79493,0 3.25,1.23122 3.25,2.75 z" ns2:ry="2.75" ns2:rx="3.25" ns2:cy="224.25" ns2:cx="449.5" id="path7444" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
              </ns0:g>
            </ns0:g>
          </ns0:g>
        </ns0:g>
        <ns0:path transform="matrix(1.0487678,0,0,1.0487678,45.282304,-29.015526)" d="m 393,646.23718 c 0,6.48935 -5.26065,11.75 -11.75,11.75 -6.48935,0 -11.75,-5.26065 -11.75,-11.75 0,-6.48934 5.26065,-11.75 11.75,-11.75 6.48935,0 11.75,5.26066 11.75,11.75 z" ns2:ry="11.75" ns2:rx="11.75" ns2:cy="646.23718" ns2:cx="381.25" id="path7446" style="color:#000000;fill:#ffffff;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:9.07692337;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
        <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.55063653;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 415.82612,622.52874 c -0.0849,0 -0.16819,1.7e-4 -0.25212,10e-4 l -0.112,0.1216 -0.16808,-0.11356 c -0.17181,0.006 -0.33805,0.0152 -0.50424,0.0272 l -0.056,0.1247 -0.21477,-0.10242 c -0.16394,0.0151 -0.32406,0.0339 -0.48089,0.0543 l 0,0.1264 -0.26146,-0.0896 c -0.15497,0.0238 -0.30674,0.0495 -0.45288,0.0784 l 0.0607,0.1247 -0.2988,-0.0752 c -0.14157,0.0317 -0.27973,0.066 -0.41087,0.10242 l 0.1168,0.1199 -0.32683,-0.0576 c -0.12555,0.0389 -0.24603,0.0801 -0.3595,0.12315 l 0.16808,0.11201 -0.35017,-0.0399 c -0.10608,0.0449 -0.20619,0.0923 -0.2988,0.14078 l 0.21943,0.10242 -0.36418,-0.0209 c -0.0843,0.0501 -0.15924,0.10213 -0.22877,0.15514 l 0.26146,0.0896 -0.36884,0 c -0.06,0.0538 -0.11454,0.10862 -0.15875,0.16474 l 0.29881,0.0736 -0.36416,0.0192 c -0.035,0.057 -0.0614,0.11384 -0.0794,0.17275 l 0.3315,0.0575 -0.35485,0.0384 c -0.004,0.0288 -0.004,0.0573 -0.004,0.0863 0,0.0291 5.2e-4,0.0575 0.004,0.0863 l 0.35485,0.0384 -0.3315,0.0575 c 0.0181,0.0588 0.0444,0.11581 0.0794,0.17273 l 0.36416,0.0192 -0.29881,0.0735 c 0.0443,0.0561 0.0987,0.11102 0.15875,0.16475 l 0.36884,0 -0.26146,0.0896 c 0.0695,0.053 0.14446,0.10509 0.22877,0.15514 l 0.36418,-0.0207 -0.21943,0.10241 c 0.0925,0.0485 0.19275,0.0958 0.2988,0.14078 l 0.35017,-0.0399 -0.16808,0.112 c 0.11342,0.043 0.234,0.0843 0.3595,0.12315 l 0.32683,-0.0576 -0.1168,0.11991 c 0.13118,0.0364 0.2693,0.0707 0.41087,0.10241 l 0.2988,-0.0752 -0.0607,0.1247 c 0.14614,0.0289 0.29791,0.0546 0.45288,0.0784 l 0.26146,-0.0896 0,0.12639 c 0.15683,0.0206 0.31695,0.0392 0.48089,0.0543 l 0.21477,-0.10241 0.056,0.12469 c 0.16619,0.0127 0.33243,0.021 0.50424,0.0272 l 0.16808,-0.11356 0.112,0.1216 c 0.0839,10e-4 0.16716,10e-4 0.25212,10e-4 0.0849,0 0.16819,-1.1e-4 0.25212,-10e-4 l 0.112,-0.1216 0.16808,0.11356 c 0.1718,-0.006 0.33805,-0.0152 0.50424,-0.0272 l 0.056,-0.12469 0.21477,0.10241 c 0.16394,-0.0151 0.32406,-0.0339 0.48089,-0.0543 l 0,-0.12639 0.26146,0.0896 c 0.15497,-0.0238 0.30673,-0.0495 0.45288,-0.0784 l -0.0607,-0.1247 0.29881,0.0752 c 0.14157,-0.0317 0.27972,-0.066 0.41086,-0.10241 l -0.11666,-0.11991 0.32682,0.0576 c 0.12554,-0.0389 0.24602,-0.0801 0.35951,-0.12315 l -0.16808,-0.112 0.35016,0.0399 c 0.10608,-0.0449 0.20619,-0.0923 0.29881,-0.14078 l -0.21943,-0.10241 0.36416,0.0207 c 0.0844,-0.0501 0.15926,-0.10199 0.22878,-0.15514 l -0.26146,-0.0896 0.36885,0 c 0.06,-0.0538 0.11454,-0.10862 0.15873,-0.16475 l -0.29881,-0.0735 0.36418,-0.0192 c 0.035,-0.057 0.0612,-0.11383 0.0794,-0.17273 l -0.3315,-0.0575 0.35485,-0.0384 c 0.004,-0.0288 0.004,-0.0573 0.004,-0.0863 0,-0.0291 -5.2e-4,-0.0575 -0.004,-0.0863 l -0.35485,-0.0384 0.3315,-0.0575 c -0.0181,-0.0588 -0.0444,-0.11581 -0.0794,-0.17275 l -0.36418,-0.0192 0.29881,-0.0736 c -0.0443,-0.0562 -0.0987,-0.11102 -0.15873,-0.16474 l -0.36885,0 0.26146,-0.0896 c -0.0695,-0.053 -0.14445,-0.10509 -0.22878,-0.15514 l -0.36416,0.0207 0.21943,-0.10241 c -0.0927,-0.0485 -0.19275,-0.0958 -0.29881,-0.14078 l -0.35016,0.0399 0.16808,-0.112 c -0.11356,-0.043 -0.23401,-0.0844 -0.35951,-0.12315 l -0.32682,0.0576 0.11666,-0.11991 c -0.13119,-0.0364 -0.26929,-0.0707 -0.41086,-0.10241 l -0.29881,0.0752 0.0607,-0.1247 c -0.14615,-0.0289 -0.29791,-0.0546 -0.45288,-0.0784 l -0.26146,0.0896 0,-0.12639 c -0.15683,-0.0206 -0.31695,-0.0392 -0.48089,-0.0543 l -0.21477,0.10241 -0.056,-0.12469 c -0.16619,-0.0127 -0.33244,-0.021 -0.50424,-0.0272 l -0.16808,0.11356 -0.112,-0.1216 c -0.0839,-0.001 -0.16714,-0.001 -0.25212,-0.001 z" id="path7448" ns1:connector-curvature="0"/>
        <ns0:path transform="matrix(-1,0,0,1,834.625,0)" ns2:open="true" ns2:end="7.609003" ns2:start="3.1415927" d="m 414.75,636.92468 c 0,-1.41523 1.14727,-2.5625 2.5625,-2.5625 1.41523,0 2.5625,1.14727 2.5625,2.5625 0,1.17585 -0.80026,2.20081 -1.941,2.48599" ns2:ry="2.5625" ns2:rx="2.5625" ns2:cy="636.92468" ns2:cx="417.3125" id="path7450" style="color:#000000;fill:#ffffff;fill-opacity:0;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      </ns0:g>
      <ns0:g style="display:inline" id="g7452" transform="matrix(0.73812401,0,0,0.73812401,380.50652,375.64387)" ns1:label="help">
        <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="cszsc" id="path7454" d="m 14.883007,5.3804864 c 0,4.5113247 -6.1837857,12.1788466 -7.884289,8.1726886 C 3.7280353,5.8478818 -1.1480278,12.785825 -3.4540023,8.2192786 -5.7318686,3.7083956 5.0017747,3.4589032 6.0524539,-0.76449404 7.5657882,-6.8476209 14.883007,0.86916191 14.883007,5.3804864 z" ns1:connector-curvature="0"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="csszz" id="path7456" d="m 49.570335,7.2077552 c 5.552326,3.1568318 -4.054237,6.3454198 -8.406364,6.3454198 -4.352128,0 -7.88429,-3.6613639 -7.88429,-8.1726886 0,-4.51132449 6.299344,-8.4568909 10.364154,-5.69282488 4.004574,2.72310568 0.30796,4.32561458 5.9265,7.52009368 z" ns1:connector-curvature="0"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="czzsc" id="path7458" d="M 14.883007,40.795492 C 10.153865,42.297569 9.5817611,52.389019 5.8507498,49.598133 1.9051658,46.646743 6.5683818,41.370391 0.39546008,42.207355 -5.749129,43.040477 -1.6161417,34.542357 6.998718,32.622802 c 4.247952,-0.946524 7.884289,3.661364 7.884289,8.17269 z" ns1:connector-curvature="0"/>
        <ns0:path style="fill:none;stroke:#000000;stroke-width:3.0788765;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" ns2:nodetypes="czzsz" id="path7460" d="m 48.695879,41.523268 c -6.690955,1.878845 -1.74186,7.467642 -6.494845,8.101936 -4.565071,0.60922 -6.451929,-4.759667 -7.063008,-8.829712 -0.607512,-4.046283 2.723221,-11.00695 6.025945,-8.17269 2.842221,2.439078 14.270309,7.008298 7.531908,8.900466 z" ns1:connector-curvature="0"/>
        <ns0:path style="fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:5.44904566;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:1.20000057" id="path7462" d="m 24.038299,-1.8893343 c -13.331156,0 -24.15066551,11.215268 -24.15066551,25.0340843 0,13.818818 10.81950951,25.034086 24.15066551,25.034086 13.331155,0 24.150665,-11.215268 24.150665,-25.034086 0,-13.8188163 -10.81951,-25.0340843 -24.150665,-25.0340843 z m 0,13.1758353 c 6.314752,-2e-6 11.439789,5.312505 11.439789,11.858249 0,6.545744 -5.125037,11.85825 -11.439789,11.85825 -6.314753,0 -11.439789,-5.312506 -11.439789,-11.85825 0,-6.545744 5.125036,-11.858249 11.439789,-11.858249 z" ns1:connector-curvature="0"/>
        <ns0:path ns2:nodetypes="ssssssssss" ns1:connector-curvature="0" d="m 24.038299,0.64151822 c -11.983426,0 -21.7091234,10.08144678 -21.7091234,22.50323178 0,12.421787 9.7256974,22.503233 21.7091234,22.503233 11.983425,0 21.709123,-10.081446 21.709123,-22.503233 0,-12.421785 -9.725698,-22.50323178 -21.709123,-22.50323178 z m 0,11.75499178 c 5.72365,-10e-7 10.368951,4.81522 10.368951,10.74824 0,5.93302 -4.645301,10.748241 -10.368951,10.748241 -5.723651,0 -10.368951,-4.815221 -10.368951,-10.748241 0,-5.93302 4.6453,-10.74824 10.368951,-10.74824 z" id="path7464" style="fill:#ffffff;fill-opacity:1;stroke:none"/>
        <ns0:path id="path7466" d="M 15.285859,2.4743562 C 10.300148,4.7510891 6.2906124,8.8924864 4.0942149,14.060578 c 4.5852109,-0.05424 7.5641511,2.312337 10.4742311,4.770797 1.039847,-2.439378 2.955558,-4.410322 5.308857,-5.488211 C 19.04958,9.2220694 17.608406,5.5277226 15.285859,2.4743562 z m 17.504879,0 c -2.236928,2.9126777 -4.141872,6.1687757 -4.591443,10.8688078 2.353298,1.077889 4.269009,3.048833 5.308856,5.488211 3.649601,-3.010131 7.184393,-4.998491 10.474231,-4.770797 C 41.785985,8.8924864 37.776449,4.7510891 32.790738,2.4743562 z M 14.568446,27.440332 c -3.491414,0.891924 -6.9828169,1.139291 -10.4742311,4.770797 2.1963975,5.16809 6.2059331,9.345358 11.1916441,11.622092 0.6226,-4.22438 1.814986,-8.080331 4.591444,-10.868809 -2.353299,-1.077889 -4.26901,-3.084703 -5.308857,-5.52408 z m 18.939705,0 c -1.039847,2.439377 -2.955558,4.446191 -5.308856,5.52408 2.320332,2.829279 3.711757,6.598889 4.591443,10.868809 4.985711,-2.276734 8.995247,-6.454002 11.191644,-11.622092 -2.4835,-2.795962 -6.191952,-4.133379 -10.474231,-4.770797 z" style="fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none" ns1:connector-curvature="0"/>
      </ns0:g>
    </ns0:g>
    <ns0:g transform="matrix(0.67009649,0,0,0.67009649,310.12555,-414.69725)" id="g7470">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:12;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path7472" ns2:cx="375.91565" ns2:cy="950.53882" ns2:rx="12.462757" ns2:ry="12.551146" d="m 388.37841,950.53882 c 0,6.9318 -5.57977,12.55114 -12.46276,12.55114 -6.88299,0 -12.46276,-5.61934 -12.46276,-12.55114 0,-6.93181 5.57977,-12.55115 12.46276,-12.55115 6.88299,0 12.46276,5.61934 12.46276,12.55115 z"/>
      <ns0:g style="display:inline" id="g7474" ns1:label="blender" transform="matrix(3.75,0,0,3.75,-789.66632,-1118.5571)">
        <ns0:path ns1:connector-curvature="0" id="path7476" transform="translate(241.0002,217)" d="m 67.8125,328.0625 c -0.24052,0.0404 -0.472023,0.15754 -0.625,0.375 -0.305953,0.43491 -0.212493,1.03265 0.21875,1.34375 l 1.6875,1.21875 -1.28125,0 -1.0625,0 -3.71875,0 C 62.473823,331 62,331.44257 62,332 c 0,0.55743 0.473823,1 1.03125,1 l 2.903109,0 -4.432138,5.08839 c -0.419418,0.48332 -0.638516,1.14294 -0.189721,1.59911 0.448795,0.45617 1.143082,0.45207 1.5625,-0.0312 l 2.4375,-2.8125 c 0.510062,1.36413 1.653338,2.50504 3.21875,2.96875 2.640781,0.78227 5.458668,-0.61365 6.28125,-3.125 0.62887,-1.91995 -0.09979,-3.93258 -1.65625,-5.125 l -4.625,-3.34375 c -0.215622,-0.15555 -0.47823,-0.19664 -0.71875,-0.15625 z m 2.1875,4 c 1.656494,0 3,1.30442 3,2.9375 0,1.63308 -1.343506,2.96875 -3,2.96875 -1.656494,0 -3,-1.33567 -3,-2.96875 0,-1.63308 1.343506,-2.9375 3,-2.9375 z" style="fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:0.5333333;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns2:nodetypes="csccccsssccsccssccccsssss"/>
        <ns0:path transform="matrix(1.8621708,0,0,1.7996949,182.32089,-49.374842)" d="m 70.023437,333.98828 c 0,0.51993 -0.416235,0.94141 -0.929687,0.94141 -0.513452,0 -0.929688,-0.42148 -0.929688,-0.94141 0,-0.51992 0.416236,-0.94141 0.929688,-0.94141 0.513452,0 0.929687,0.42149 0.929687,0.94141 z" ns2:ry="0.94140625" ns2:rx="0.9296875" ns2:cy="333.98828" ns2:cx="69.09375" id="path7478" style="fill:#000000;fill-opacity:1;stroke:none" ns2:type="arc"/>
      </ns0:g>
    </ns0:g>
    <ns0:g ns1:label="file-roller" transform="matrix(0.67009649,0,0,0.67009649,310.3109,-385.36407)" id="g7480">
      <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 346.83588,794.44498 -4.77297,15.55635 c 0.18303,3.76817 1.70957,7.45731 4.24264,10.25305 3.07474,3.39357 7.61825,5.40802 12.19759,5.40802 4.57934,0 9.12285,-2.01445 12.19759,-5.40802 l -0.88388,-14.31891 6.71751,-12.72792 -29.69848,1.23743" id="path7482" ns1:path-effect="#path-effect30843" ns1:original-d="m 346.83588,794.44498 -4.77297,15.55635 c 0,0 3.53553,10.78338 4.24264,10.25305 0.7071,-0.53033 24.39518,0 24.39518,0 l -0.88388,-14.31891 6.71751,-12.72792 z" ns1:connector-curvature="0"/>
      <ns0:g transform="matrix(3.9852721,0,0,3.9852721,-950.24365,71.174473)" style="display:inline" id="g7484" ns1:label="file-roller">
        <ns0:rect transform="translate(241.0002,217)" y="-42" x="82" height="16" width="16" id="rect7486" style="fill:none;stroke:none"/>
        <ns0:path ns1:r_cy="true" ns1:r_cx="true" ns2:nodetypes="czcszccccccc" id="path7488" d="m 330.07659,187.00703 c 0,0 -2.91924,-0.0221 -3.10498,-0.0221 -0.18574,0 -0.26784,0.0324 -0.37159,-0.14741 -0.30689,-0.42982 -0.52143,-1.10364 -0.57752,-1.71708 -0.0109,-0.11882 -0.20696,-0.12631 -0.30151,-0.12683 L 323.15958,185 c -0.13341,0 -0.15695,0.24121 -0.15695,0.24121 -0.0519,1.89982 0.71945,4.7556 2.88858,4.74728 L 333.7812,190 c -2.67921,-0.16112 -2.63112,-1.34814 -2.84212,-2.47213 -0.18112,-0.35221 -0.25941,-0.52078 -0.5697,-0.52078 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none;stroke-width:0.62873191;marker:none;visibility:visible;display:inline;overflow:visible" ns1:connector-curvature="0"/>
        <ns0:path style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" d="m 332.0002,181.49621 2.5,0 c 3.80719,0 4.21897,8 0,8 l -2.9375,0" id="path7490" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
        <ns0:path ns2:nodetypes="csscccsccccsccccccsc" ns1:connector-curvature="0" id="path7492" transform="translate(241.0002,217)" d="m 85.09375,-36 c -1.27743,0 -2.3125,2.02507 -2.3125,4.5 0,2.47494 1.03507,4.375 2.3125,4.375 0.0306,0 0.06355,-0.02925 0.09375,-0.03125 l 0,0.03125 8.812498,-0.875 c -1.8125,0 -3.062498,-1.098645 -3.062498,-3.5 0,-2.389424 1.03608,-3.5 3.062498,-3.5 l -1.585934,-0.996098 C 89.184425,-36.006039 85.09375,-36 85.09375,-36 z m 0.02344,0.992187 4.97656,0.0078 c 0.16968,2.66e-4 0.32247,0.18898 0.1875,0.375 -0.84239,1.515638 -0.897612,3.781759 -0.356694,5.569432 0,0.17445 -0.14283,0.3125 -0.3125,0.3125 l -5.048906,0.01386 c -0.16969,0 -0.25,-0.20055 -0.25,-0.375 -0.0858,-1.75606 -0.921312,-4.157719 0.585288,-5.841109 0,0 0.04901,-0.06277 0.218752,-0.0625 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.34051171;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
        <ns0:path ns2:nodetypes="cccccccccccccccccccsccc" id="path7494" d="m 330.00832,177 c -0.39473,0 -0.70961,0.17025 -0.88958,0.46259 l -2.28241,3.68924 -0.14046,0.27756 0.30433,0 1.10135,0 0.11704,0 0.0469,-0.10414 1.4538,-2.17057 c 0.0363,-0.0581 0.15888,-0.15034 0.28091,-0.15034 l 7.3961,0.003 c 0.0786,-0.005 0.079,0.10987 0.079,0.10987 l -2.87252,5.72088 -0.0937,0.16191 0.16385,0.0926 0.0698,0.70127 0.6942,0.36803 0.0936,-0.1619 3.46967,-7 c 0.13852,-0.23162 0.005,-1.3902 -0.10814,-1.59514 -0.12605,-0.22734 -0.3837,-0.41187 -0.71398,-0.40478 l -8.16989,0 z" style="fill:#000000;fill-opacity:1;fill-rule:evenodd;stroke:none" ns1:connector-curvature="0"/>
        <ns0:path d="M 35.5625,31.953125 C 35.5625,33.635868 34.765007,35 33.78125,35 32.797493,35 32,33.635868 32,31.953125 c 0,-1.682743 0.797493,-3.046875 1.78125,-3.046875 0.983757,0 1.78125,1.364132 1.78125,3.046875 z" ns2:ry="3.046875" ns2:rx="1.78125" ns2:cy="31.953125" ns2:cx="33.78125" id="path7496" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc" transform="matrix(0.49627604,0,0,0.49230822,318.11937,169.76921)"/>
      </ns0:g>
    </ns0:g>
    <ns0:g transform="matrix(3.9991698,0,0,3.9991698,92.8635,350.39362)" ns1:label="#g5607" id="default-pointer-c-1" style="display:inline" ns1:export-filename="/home/jimmac/gfx/redhat/redhat-ux/Products/RHEL/RHEL7/video-jingles/tex/pointer.png" ns1:export-xdpi="90" ns1:export-ydpi="90">
      <ns0:path style="color:#000000;fill:url(#linearGradient14910-9);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path5565-2" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
      <ns0:path ns2:nodetypes="cccccccc" id="path6242-4" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:g ns1:export-ydpi="90" ns1:export-xdpi="90" transform="translate(499,-725)" style="display:inline" id="vpn" ns1:label="network-vpn">
      <ns0:g style="fill:#bebebe;fill-opacity:1" transform="translate(181,233)" ns1:label="lock" id="g13201">
        <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" id="rect13203" width="16" height="16" x="20" y="276" ns1:label="a"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="cc" ns1:connector-curvature="0" id="path12679-6" d="m 208.99975,519 0,3" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible"/>
      <ns0:path ns1:connector-curvature="0" id="path12681-3" d="m 202.99975,523 12,0" style="color:#bebebe;fill:none;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible"/>
      <ns0:rect ry="0" transform="translate(-2.5e-4,272)" y="242" x="205" height="6" width="8" id="rect13312" style="color:#bebebe;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible"/>
      <ns0:path style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#bebebe;fill:#000000;fill-opacity:1;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans" d="m 208.99977,510.00041 c -1.64501,0 -3,1.355 -3,3 l 0,2 0,1.00001 1,0 4,0 1,0 0,-1.00001 0,-2 c 0,-1.645 -1.35499,-3 -3,-3 z m 0,2 c 0.56413,0 1,0.43588 1,1 l 0,1 -2,0 0,-1 c 0,-0.56412 0.43587,-1 1,-1 z" id="path13314" ns1:connector-curvature="0"/>
    </ns0:g>
    <ns0:g id="g12006">
      <ns0:g id="g5525" transform="translate(689,-168)" ns1:label="audio-volume-medium" style="display:inline">
        <ns0:path ns2:nodetypes="ccccccccc" id="path5533" d="m 20,222 2.484375,0 2.968754,-3 0.546871,0.0156 0,11 -0.475297,8.3e-4 L 22.484375,227 20,227 l 0,-5 z" style="color:#bebebe;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" ns1:connector-curvature="0"/>
        <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" id="rect5535" width="16" height="16" x="20" y="217" ns1:label="audio-volume-high"/>
        <ns0:path clip-path="url(#clipPath6279-7-9)" ns2:type="arc" style="fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path3718-5" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
        <ns0:path clip-path="url(#clipPath6265-3-4)" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3726-1" style="fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" ns2:type="arc" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
        <ns0:path clip-path="url(#clipPath6259-8-81)" ns2:type="arc" style="opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path3728-0" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
      </ns0:g>
      <ns0:g transform="translate(689,-639)" ns1:label="system-shutdown" id="g4692-3" style="display:inline">
        <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect10837-3-0" y="688" x="40" ry="0.15129246" rx="0.14408804" height="16" width="16"/>
        <ns0:path ns2:open="true" ns2:end="10.471045" ns2:start="5.239857" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" d="m 51.52343,689.95141 c 3.340544,1.94594 4.471097,6.23148 2.52516,9.57202 -1.945936,3.34054 -6.231476,4.4711 -9.57202,2.52516 -3.340544,-1.94594 -4.471097,-6.23148 -2.52516,-9.57202 0.612757,-1.05191 1.489249,-1.92583 2.542951,-2.53549" ns2:ry="7" ns2:rx="7" ns2:cy="696" ns2:cx="48" id="path3869-2" style="color:#000000;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
        <ns0:path ns2:nodetypes="cc" id="path4710" d="m 48,689 0,5" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:g id="g12661" transform="translate(666.07286,-166.91767)" ns1:label="network-wired" style="display:inline">
        <ns0:rect ns1:label="audio-volume-high" y="217" x="20" height="16" width="16" id="rect12673" style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible"/>
        <ns0:path id="rect12675" transform="translate(80,257)" d="m -55.25,-40 c -0.952203,0 -1.75,0.7978 -1.75,1.75 l 0,4.5 c 0,0.9522 0.797797,1.75 1.75,1.75 l 0.125,0 -0.78125,1.5625 -0.71875,1.4375 1.625,0 6,0 1.625,0 -0.71875,-1.4375 L -48.875,-32 l 0.125,0 c 0.952203,0 1.75,-0.7978 1.75,-1.75 l 0,-4.5 c 0,-0.9522 -0.797797,-1.75 -1.75,-1.75 l -6.5,0 z m 0.25,2 6,0 0,4 -6,0 0,-4 z" style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#bebebe;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans" ns1:connector-curvature="0"/>
        <ns0:path style="color:#bebebe;fill:none;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible" d="m 88,196 0,4" id="path12679" transform="translate(-60.0003,30)" ns1:connector-curvature="0"/>
        <ns0:path style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible" d="m 21.99975,231 12,0" id="path12681" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="rect12003" d="m 759.10724,57.4163 -3.74999,3.750004 -3.75001,-3.750005 z" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:g>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer5" ns1:label="play" ns2:insensitive="true" style="display:inline">
    <ns0:g style="display:inline" transform="matrix(2.862069,0,0,2.862069,49.362076,-2561.8469)" id="g4607">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:0.74427478;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path2086" ns2:cx="122" ns2:cy="79" ns2:rx="29" ns2:ry="29" d="m 151,79 c 0,16.016258 -12.98374,29 -29,29 -16.01626,0 -29,-12.983742 -29,-29 0,-16.016258 12.98374,-29 29,-29 16.01626,0 29,12.983742 29,29 z" transform="translate(7.5,897.86218)"/>
      <ns0:g transform="matrix(2.46875,0,0,2.46875,13.25,-244.41907)" ns1:label="media-playback-start" id="g4135" style="display:inline">
        <ns0:path style="font-size:xx-small;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Bitstream Vera Sans;-inkscape-font-specification:Bitstream Vera Sans" d="m 84,609 0,10 0.90625,0 L 85,619 c 0.174914,10e-4 0.347782,-0.0388 0.5,-0.125 l 7,-4 c 0.310699,-0.17189 0.46875,-0.52345 0.46875,-0.875 0,-0.35155 -0.158051,-0.70311 -0.46875,-0.875 l -7,-4 C 85.347782,609.03875 85.174914,608.99869 85,609 l -0.09375,0 z" transform="translate(-39.99995,-119)" id="path3807-1-1-9-38-4" ns1:connector-curvature="0" ns2:nodetypes="ccccccsccccc"/>
      </ns0:g>
    </ns0:g>
  </ns0:g>
</ns0:svg>
