<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Nätkonton</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Nätkonton</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan mata in dina kontouppgifter för vissa nättjänster, så som Google och Facebook, i fönstret <span class="app">Nätkonton</span>. Detta kommer att låta dig använda program för att nå nättjänster som e-post, kalendrar, chatt och dokument.</p>
<div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="accounts-add.html" title="Lägg till ett konto"><span class="title">Lägg till ett konto</span><span class="linkdiv-dash"> — </span><span class="desc">Tillåt program att få åtkomst till dina nätkonton för foton, kontakter, kalendrar och så vidare.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="accounts-remove.html" title="Ta bort ett konto"><span class="title">Ta bort ett konto</span><span class="linkdiv-dash"> — </span><span class="desc">Ta bort tillgång till en nättjänstleverantör från dina program.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="accounts-whyadd.html" title="Varför lägga till ett konto?"><span class="title">Varför lägga till ett konto?</span><span class="linkdiv-dash"> — </span><span class="desc">Varför ska jag lägga till e-post eller sociala media-konton i min skrivbordsmiljö?</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="accounts-which-application.html" title="Nättjänster och program"><span class="title">Nättjänster och program</span><span class="linkdiv-dash"> — </span><span class="desc">Program kan använda de konton som skapats i <span class="app">Nätkonton</span> och tjänsterna de utnyttjar.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="accounts-disable-service.html" title="Styr vilka nättjänster ett konto kan användas med"><span class="title">Styr vilka nättjänster ett konto kan användas med</span><span class="linkdiv-dash"> — </span><span class="desc">Vissa nätkonton kan användas för att nå flera tjänster (exempelvis kalender och e-post). Du kan styra vilken av dessa tjänster som kan användas av program.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="accounts-provider-not-available.html" title="Varför är min kontotyp inte på listan?"><span class="title">Varför är min kontotyp inte på listan?</span><span class="linkdiv-dash"> — </span><span class="desc">Vad gör jag om en nättjänsteleverantör inte finns på listan?</span></a></div>
</div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html" title="Användarkonton">användarkonton</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="net-chat.html" title="Chatt &amp; sociala medier">Chatt &amp; sociala medier</a><span class="desc"> — 
      <span class="link"><a href="net-chat-empathy.html" title="Snabbmeddelanden på Ubuntu">Chat on any network using <span class="app">Empathy</span></a></span>,
      <span class="link"><a href="net-chat-video.html" title="Videosamtal">make video calls</a></span>,
      <span class="link"><a href="net-chat-skype.html" title="Hur använder jag Skype på Ubuntu?">install skype</a></span>
    </span>
</li>
<li class="links "><a href="gs-connect-online-accounts.html" title="Ansluta till nätkonton">En handledning i att ansluta till nätkonton</a></li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
