<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Dela ditt skrivbord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="prefs-sharing.html.sv" title="Dela-inställningar">Dela-inställningar</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a> » <a class="trail" href="sharing.html.sv" title="Dela">Dela</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Dela ditt skrivbord</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan låta andra personer se och styra ditt skrivbord från en annan dator med ett skrivbordsvisningsprogram. Konfigurera <span class="gui">Skärmdelning</span> till att låta andra personer få åtkomst till ditt skrivbord och ställ in säkerhetsinställningarna.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Du måste ha paketet <span class="app">Vino</span> installerat för att <span class="gui">Skärmdelning</span> ska visas.</p></div></div></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Dela</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Dela</span> för att öppna panelen.</p></li>
<li class="steps">
<p class="p">Om <span class="gui">Dela</span> är <span class="gui">AV</span>, slå om den till <span class="gui">PÅ</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om texten nedanför <span class="gui">Datornamn</span> låter dig redigera den, kan du <span class="link"><a href="sharing-displayname.html.sv" title="Ställ in visningsnamnet för din dator">ändra</a></span> namnet din dator visar på nätverket.</p></div></div></div></div>
</li>
<li class="steps"><p class="p">Välj <span class="gui">Skärmdelning</span>.</p></li>
<li class="steps"><p class="p">För att låta andra se ditt skrivbord, slå om <span class="gui">Skärmdelning</span> till <span class="gui">PÅ</span>. Detta innebär att andra personer kan försöka att ansluta till din dator och se vad som finns på din skärm.</p></li>
<li class="steps">
<p class="p">För att låta andra interagera med ditt skrivbord, slå om <span class="gui">Tillåt fjärrkontroll</span> till <span class="gui">PÅ</span>. Detta låter den andra personen att flytta din mus, köra program och bläddra bland filer på din dator, beroende på säkerhetsinställningarna som du använder för närvarande.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Detta alternativ är aktiverat som standard när <span class="gui">Skärmdelning</span> är <span class="gui">PÅ</span>.</p></div></div></div></div>
</li>
</ol></div></div></div>
</div>
<div id="security" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Säkerhet</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Det är viktigt att du funderar på den fulla vidden av vad varje säkerhetsalternativ innebär innan du ändrar det.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Nya anslutningar måste be om åtkomst</dt>
<dd class="terms">
<p class="p">Om du vill kunna välja huruvida någon ska beviljas åtkomst till ditt skrivbord, aktivera <span class="gui">Nya anslutningar måste fråga efter åtkomst</span>. Om du inaktiverar detta alternativ kommer du inte att blir tillfrågad huruvida du vill tillåta någon att ansluta till din dator.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Detta alternativ är aktiverat som standard.</p></div></div></div></div>
</dd>
<dt class="terms">Kräv ett lösenord</dt>
<dd class="terms">
<p class="p">För att kräva att andra personer använder ett lösenord när de ansluter till ditt skrivbord, aktivera <span class="gui">Begär lösenord</span>. Om du inte använder detta alternativ kan vem som helst försöka se ditt skrivbord.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Detta alternativ är inaktiverat som standard, men du bör aktivera det och ställa in ett säkert lösenord.</p></div></div></div></div>
</dd>
</dl></div></div></div>
</div></div>
</div></div>
<div id="networks" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Nätverk</span></h2></div>
<div class="region"><div class="contents"><p class="p">Sektionslistan <span class="gui">Nätverk</span> listar nätverken som du för närvarande är ansluten till. Använd <span class="gui">ON | OFF</span>-knappen intill respektive för att välja var ditt skrivbord kan delas.</p></div></div>
</div></div>
<div id="notification-icon" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Sluta dela ditt skrivbord</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan koppla från någon som ser ditt skrivbord via <span class="gui">aviseringsikonen</span> i meddelandefältet. För att göra detta:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna meddelandefältet genom att trycka <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>M</kbd></span></span>, eller genom att flytta din musmarkör längst ner på skärmen.</p></li>
<li class="steps"><p class="p">Klicka på ikonen <span class="gui">Skrivbord</span> i <span class="gui">meddelandefältet</span>. Detta öppnar panelen <span class="app">Dela</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Skärmdelning</span>.</p></li>
<li class="steps"><p class="p">Slå om skjutreglaget <span class="gui">Skärmdelning</span> till <span class="gui">AV</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="sharing.html.sv" title="Dela">Dela</a><span class="desc"> — <span class="link"><a href="sharing-desktop.html.sv" title="Dela ditt skrivbord">Skrivbordsdelning</a></span>, <span class="link"><a href="files-share.html.sv" title="Dela filer visa e-post">Dela filer via e-post</a></span>, <span class="link"><a href="sharing-media.html.sv" title="Dela din musik, foton och videor">Mediadelning</a></span>…</span>
</li>
<li class="links ">
<a href="prefs-sharing.html.sv" title="Dela-inställningar">Dela-inställningar</a><span class="desc"> — <span class="link"><a href="sharing-bluetooth.html.sv" title="Styr delning över Bluetooth">Bluetooth-delning</a></span>, <span class="link"><a href="sharing-personal.html.sv" title="Dela ut dina personliga filer">Delning av personliga filer</a></span>, <span class="link"><a href="sharing-desktop.html.sv" title="Dela ditt skrivbord">Skärmdelning</a></span>, <span class="link"><a href="sharing-media.html.sv" title="Dela din musik, foton och videor">Mediadelning</a></span>…</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
