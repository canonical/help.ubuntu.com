<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Instruktioner för att para ihop specifika enheter</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 23.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="bluetooth.html.sv" title="Bluetooth">Bluetooth</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Instruktioner för att para ihop specifika enheter</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Även om du lyckas hitta manualen för enheten är det inte säkert att den innehåller tillräckligt med information för att genomföra en framgångsrik ihopparning. Här kommer detaljer för ett antal vanliga enheter.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">PlayStation 5-handkontroller</dt>
<dd class="terms"><p class="p">Håll ner <span class="media"><span class="media media-image"><img src="figures/ps-create.svg" class="media media-inline" alt="Create"></span></span>-knappen och tryck på <span class="media"><span class="media media-image"><img src="figures/ps-button.svg" class="media media-inline" alt="PS"></span></span>-knappen tills ljuspanelen blinkar för att göra den synlig och para ihop den som vilken annan Bluetooth-enhet som helst.</p></dd>
<dt class="terms">PlayStation 4-handkontroller</dt>
<dd class="terms">
<p class="p">Kombinationen av <span class="media"><span class="media media-image"><img src="figures/ps-button.svg" class="media media-inline" alt="PS"></span></span>- och ”Share”-knapparna för att para ihop handkontrollen kan också användas för att göra handkontrollen synlig och para ihop den som vilken annan Bluetooth-enhet som helst.</p>
<p class="p">De enheterna kan också använda ”kabel-ihopparning”. Anslut handkontrollerna via USB med <span class="gui">Bluetoothinställningar</span> öppnat och Bluetooth påslaget. Du kommer att tillfrågas huruvida du vill installera handkontrollerna utan att behöva trycka på <span class="media"><span class="media media-image"><img src="figures/ps-button.svg" class="media media-inline" alt="PS"></span></span>-knappen. Koppla från dem och tryck på <span class="media"><span class="media media-image"><img src="figures/ps-button.svg" class="media media-inline" alt="PS"></span></span>-knappen för att använda dem över Bluetooth.</p>
</dd>
<dt class="terms">PlayStation 3-handkontroller</dt>
<dd class="terms"><p class="p">De enheterna använder ”kabel-ihopparning”. Anslut handkontrollerna via USB med <span class="gui">Bluetoothinställningar</span> öppnat och Bluetooth påslaget. Efter att ha tryckt på <span class="media"><span class="media media-image"><img src="figures/ps-button.svg" class="media media-inline" alt="PS"></span></span>-knappen kommer du att tillfrågas huruvida du vill installera handkontrollerna. Koppla från dem och tryck på <span class="media"><span class="media media-image"><img src="figures/ps-button.svg" class="media media-inline" alt="PS"></span></span>-knappen för att använda dem över Bluetooth.</p></dd>
<dt class="terms">PlayStation 3 BD-fjärrkontroll</dt>
<dd class="terms"><p class="p">Håll ner ”Start”- och ”Enter”-knapparna samtidigt under cirka fem sekunder. Du kan sen välja fjärrkontrollen i enhetslistan som vanligt.</p></dd>
<dt class="terms">Nintendo Wii- och Wii U-fjärrkontroller</dt>
<dd class="terms"><p class="p">Använd den röda ”Sync”-knappen bakom batteriluckan för att starta ihopparningsprocessen. Andra knappkombinationer kommer inte att behålla ihopparningsinformationen så du skulle komma att behöva att göra om det igen inom kort. Notera också att viss programvara som konsolemulatorer vill ha direktåtkomst till fjärrkontrollerna, och i de fallen bör du inte installera dem direkt i Bluetooth-panelen. Referera till programmets handbok för instruktioner.</p></dd>
<dt class="terms">ION iCade</dt>
<dd class="terms"><p class="p">Håll nere de nedre fyra knapparna och den övre vita knappen för att starta ihopparningsprocessen. Se till att när ihopparningsinstruktionerna visas bara använda kardinalriktningarna för att mata in koden, följt av någon av de två vita knapparna längst till höger om arkadspaken för att bekräfta.</p></dd>
</dl></div></div></div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="bluetooth.html.sv" title="Bluetooth">Bluetooth</a><span class="desc"> — Anslut till enheter över Bluetooth för att överföra filer eller använda trådlöst ljud.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="bluetooth-visibility.html.sv" title="Vad är Bluetooth-synlighet?">Vad är Bluetooth-synlighet?</a><span class="desc"> — Huruvida andra enheter kan detektera din dator.</span>
</li></ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
