<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Resurser</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = "index.html.en";
        } else {
                window.location = href.replace(/\.html.*/, ".html.en");
        }
         return false;
      }
      function browserPreferredLanguage() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = href;
        } else {
                window.location = href.replace(/\.html.*/, ".html");
        }
        return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../18.04" class="trail">Ubuntu 18.04</a> » <a class="trail" href="index.html.sv" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="cgroups.html.sv" title="Control Groups">Control Groups</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups-manager.html.sv" title="Manager">Föregående</a><a class="nextlinks-next" href="clustering.html.sv" title="Kluster">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Resurser</h1></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
          <p class="para">Manual pages referenced above can be found at:</p>
          <div class="screen"><pre class="contents "><a href="http://manpages.ubuntu.com/manpages/en/man8/cgm.1.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/cgm.1.html">cgm</a>
<a href="http://manpages.ubuntu.com/manpages/en/man5/cgconfig.conf.5.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man5/cgconfig.conf.5.html">cgconfig.conf</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/cgmanager.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/cgmanager.8.html">cgmanager</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/cgproxy.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/cgproxy.8.html">cgproxy</a>
</pre></div>
        </li>
<li class="list itemizedlist">
          <p class="para">The upstream cgmanager project is hosted at <a href="http://cgmanager.linuxcontainers.org" class="ulink" title="http://cgmanager.linuxcontainers.org">linuxcontainers.org</a>.</p>
        </li>
<li class="list itemizedlist">
          <p class="para">The upstream kernel documentation page on cgroups can be seen <a href="https://git.kernel.org/cgit/linux/kernel/git/torvalds/linux.git/tree/Documentation/cgroups" class="ulink" title="https://git.kernel.org/cgit/linux/kernel/git/torvalds/linux.git/tree/Documentation/cgroups">here
	  </a>.</p>
        </li>
<li class="list itemizedlist">
          <p class="para">The freedesktop.org control group usage guidelines can be seen <a href="http://www.freedesktop.org/wiki/Software/systemd/PaxControlGroups/" class="ulink" title="http://www.freedesktop.org/wiki/Software/systemd/PaxControlGroups/">here</a>.</p>
        </li>
</ul></div></div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups-manager.html.sv" title="Manager">Föregående</a><a class="nextlinks-next" href="clustering.html.sv" title="Kluster">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address
          so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>
          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p>
</div>
</div>
</body>
</html>
