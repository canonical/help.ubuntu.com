<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Visa andra tidszoner</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="clock.html" title="Datum &amp; tid">Datum &amp; tid</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Visa andra tidszoner</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du vill veta vad klockan är i olika städer världen över kan du lägga till ytterligare tidszoner till klockmenyn. Dessa extrastäder kommer visas nedanför kalendern när du klickar på klockan.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på klockan och välj <span class="gui">Datum- &amp; tidsinställningar</span>.</p></li>
<li class="steps"><p class="p">Gå till fliken <span class="gui">Klocka</span> och välj <span class="gui">Tid på andra platser</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Välj platser</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">+</span> för att lägga till en plats.</p></li>
<li class="steps"><p class="p">Fyll i Platsfältet med namnet på staden du vill lägga till. Vänta en stund på att listan över möjliga träffar visas i den utfällbara listan.</p></li>
<li class="steps"><p class="p">Välj staden du vill ha, så fylls tiden på den platsen i automatiskt.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">-</span> för att ta bort en stad från listan.</p></li>
<li class="steps"><p class="p">Du kan också dra-och-släppa städerna i det här <span class="gui">Platsfönstret</span> för att ändra ordningen de visas i på klockmenyn.</p></li>
</ol></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="clock.html" title="Datum &amp; tid">Datum &amp; tid</a><span class="desc"> — <span class="link"><a href="clock-set.html" title="Ändra tid och datum">Ange datum och tid</a></span>, <span class="link"><a href="clock-timezone.html" title="Visa andra tidszoner">tidszon</a></span>, <span class="link"><a href="clock-calendar.html" title="Kalendermöten">kalender och möten</a></span>...</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="clock-set.html" title="Ändra tid och datum">Ändra tid och datum</a><span class="desc"> — Uppdatera tid/datum som visas överst i skärmen.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
