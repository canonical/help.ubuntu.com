<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" height="500" id="svg10075" version="1.1" width="840" ns2:docname="gs-datetime.svg" ns1:version="0.92.4 5da689c313, 2019-01-14">
  <ns0:defs id="defs10077">
    <ns0:linearGradient id="RHEL7" ns3:paint="gradient">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop id="stop11074" offset="0" style="stop-color:#eeedec;stop-opacity:1;"/>
      <ns0:stop id="stop11076" offset="1" style="stop-color:#eeedec;stop-opacity:1"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop id="stop7012" offset="0" style="stop-color:#eeedec;stop-opacity:0;"/>
      <ns0:stop id="stop7014" offset="1" style="stop-color:#eeedec;stop-opacity:0"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" gradientUnits="userSpaceOnUse" id="linearGradient7064" x1="-18.33782" x2="713.42853" y1="490.54935" y2="490.54935" ns1:collect="always" ns4:href="#GNOME"/>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient5885" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop id="stop5718" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17441" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop id="stop17445" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop17447" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17453" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17455" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:filter color-interpolation-filters="sRGB" height="1.1308649" id="filter5601" width="1.2058235" x="-0.10291173" y="-0.065432459" ns1:collect="always">
      <ns0:feGaussianBlur id="feGaussianBlur5603" stdDeviation="0.610872" ns1:collect="always"/>
    </ns0:filter>
    <ns0:linearGradient gradientTransform="matrix(1.0281734,0,0,1.0281734,637.14345,666.93836)" gradientUnits="userSpaceOnUse" id="linearGradient17453-7" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716-4"/>
    <ns0:linearGradient id="linearGradient5716-4">
      <ns0:stop id="stop5718-1" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720-6" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(1.0281734,0,0,1.0281734,637.14345,666.93836)" gradientUnits="userSpaceOnUse" id="linearGradient17455-1" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716-4"/>
    <ns0:linearGradient id="linearGradient16929">
      <ns0:stop id="stop16931" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop16933" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
  </ns0:defs>
  <ns2:namedview bordercolor="#666666" borderlayer="true" borderopacity="1.0" fit-margin-bottom="0" fit-margin-left="0" fit-margin-right="0" fit-margin-top="0" height="0px" id="base" pagecolor="#eeeeec" showgrid="false" width="0px" ns1:current-layer="g4890" ns1:cx="154.72357" ns1:cy="347.41188" ns1:document-units="px" ns1:pageopacity="1" ns1:pageshadow="2" ns1:showpageshadow="false" ns1:window-height="1403" ns1:window-maximized="1" ns1:window-width="2560" ns1:window-x="2560" ns1:window-y="0" ns1:zoom="1">
    <ns1:grid empspacing="5" enabled="true" id="grid17504" snapvisiblegridlinesonly="true" type="xygrid" visible="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true" ns1:groupmode="layer" ns1:label="bg">
    <ns0:rect height="656" id="background" style="fill:url(#BLANK);" width="866" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g id="layer2" transform="translate(0,-540)" ns1:groupmode="layer" ns1:label="fg">
    <ns0:g id="g11020" transform="translate(-89,-139.36217)">
      <ns0:circle cx="120" cy="278" id="path11014" r="17" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;enable-background:accumulate" transform="translate(2,453.36217)"/>
      <ns0:text id="text11016" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" xml:space="preserve"><ns0:tspan id="tspan11018" style="font-size:14px;line-height:1.25" x="122.29289" y="736.36218" ns2:role="line">3</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g id="g4890" style="display:inline" transform="matrix(2.6833333,0,0,2.6833333,-1275.5101,-1072.8539)">
      <ns0:path d="m 506.43234,611.75299 h 258.32299 c 2.21601,0 4,1.784 4,4 v 161.22982 h -4 -258.32299 -4 V 615.75299 c 0,-2.216 1.784,-4 4,-4 z" id="path5430" style="display:inline;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-opacity:1" ns2:nodetypes="sssccccss" ns1:connector-curvature="0"/>
      <ns0:path d="M 502.98343,630.36169 H 768.47408" id="path5361" style="display:inline;fill:none;stroke:#000000;stroke-width:1.01455009;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
      <ns0:path d="m 756.48074,617.84776 h 0.74998 c 0.008,-9e-5 0.0156,-3.5e-4 0.0234,0 0.19121,0.008 0.38239,0.0964 0.51561,0.23437 l 1.71089,1.71088 1.73432,-1.71088 c 0.19921,-0.17287 0.335,-0.22912 0.51561,-0.23437 h 0.74998 v 0.74998 c 0,0.21484 -0.0258,0.41297 -0.1875,0.56248 l -1.71088,1.71089 1.68745,1.68745 c 0.14113,0.14112 0.21092,0.34008 0.21093,0.53905 v 0.74997 h -0.74998 c -0.19897,0 -0.39793,-0.0698 -0.53905,-0.21093 l -1.71088,-1.71089 -1.71089,1.71089 c -0.14112,0.14114 -0.34009,0.21093 -0.53905,0.21093 h -0.74998 v -0.74997 c 0,-0.19897 0.0698,-0.39793 0.21094,-0.53905 l 1.71088,-1.68745 -1.71088,-1.71089 c -0.15806,-0.14597 -0.22737,-0.35193 -0.21094,-0.56248 z" id="path5375" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.3358984;marker:none;enable-background:new" ns2:nodetypes="ccccccccscccccscccscsccccc" ns1:connector-curvature="0"/>
      <ns0:text id="text12012" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="669.13416" y="622.67847" xml:space="preserve"><ns0:tspan id="tspan12014" style="font-size:5.21739101px;line-height:1.25" x="669.13416" y="622.67847" ns2:role="line">Datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:rect height="93.540375" id="rect9293" rx="0" ry="0" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.7453416;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" width="147.9503" x="600.56281" y="634.97662"/>
      <ns0:text id="text26176" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="645.52429" xml:space="preserve"><ns0:tspan id="tspan26178" style="font-size:5.21739101px;line-height:1.25" x="610.1059" y="645.52429" ns2:role="line">Automatisk datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:text id="text26182" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#babdb6;fill-opacity:1;stroke:none" x="610.1059" y="652.2323" xml:space="preserve"><ns0:tspan id="tspan26184" style="font-size:4.47205019px;line-height:1.25" x="610.1059" y="652.2323" ns2:role="line">Kräver internetåtkomst</ns0:tspan></ns0:text>
      <ns0:g id="g9286" transform="translate(-17.515526,-52.919256)">
        <ns0:g id="g3921" style="display:inline" transform="matrix(0.37267081,0,0,0.37267081,493.07637,552.48134)"/>
      </ns0:g>
      <ns0:rect height="5.9627328" id="rect10837-5-8-1" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.3726708;marker:none;enable-background:new" transform="scale(-1,1)" width="5.9627328" x="-514.0741" y="617.82538"/>
      <ns0:path d="m 512.58846,618.5707 h -0.37267 c -0.004,-4e-5 -0.008,-1.7e-4 -0.0117,0 -0.095,0.004 -0.19001,0.0479 -0.25621,0.11646 l -2.34696,2.13121 2.34698,2.13121 c 0.0701,0.0701 0.16899,0.10482 0.26786,0.10482 h 0.37267 v -0.37267 c 0,-0.0989 -0.0347,-0.19774 -0.10481,-0.26786 l -1.79962,-1.5955 1.79962,-1.59549 c 0.0785,-0.0725 0.11297,-0.17488 0.10481,-0.27951 z" id="path10839-9-9-5" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.66381985;marker:none;enable-background:new" ns2:nodetypes="ccsccccccccccc" ns1:connector-curvature="0"/>
      <ns0:rect height="11.925466" id="rect15386" rx="1.4906832" ry="1.4906832" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.3726708;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" width="11.925466" x="505.35666" y="615.02734"/>
      <ns0:path d="M 600.56278,658.59462 H 748.51309" id="path9309" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
      <ns0:text id="text9311" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="667.88458" xml:space="preserve"><ns0:tspan id="tspan9313" style="font-size:5.21739101px;line-height:1.25" x="610.1059" y="667.88458" ns2:role="line">Automatisk tidszon</ns0:tspan></ns0:text>
      <ns0:text id="text9315" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#babdb6;fill-opacity:1;stroke:none" x="610.1059" y="674.59259" xml:space="preserve"><ns0:tspan id="tspan9317" style="font-size:4.47205019px;line-height:1.25" x="610.1059" y="674.59259" ns2:role="line">Kräver internetåtkomst</ns0:tspan></ns0:text>
      <ns0:path d="M 600.56278,680.95488 H 748.51309" id="path9331" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
      <ns0:rect height="10.92049" id="rect939" rx="5.4602423" ry="5.4602423" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" width="19.803892" x="719.65601" y="665.09509"/>
      <ns0:circle cx="733.60791" cy="670.55194" id="circle941" r="4.4139271" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:path d="M 97.089832,2.8483222 V 19.288556 l 3.712308,-3.623922 2.12132,4.331029 c 0.5196,1.171377 3.22086,0.229524 2.45278,-1.336875 l -2.09922,-4.496756 h 4.68458 z" id="path5567" style="color:#000000;display:block;overflow:visible;visibility:visible;opacity:0.6;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;filter:url(#filter5601);enable-background:accumulate" transform="matrix(1.0281734,0,0,1.0281734,637.14345,666.93836)" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
      <ns0:path d="m 736.42336,669.32166 v 16.90341 l 3.8169,-3.72602 2.18109,4.45305 c 0.53423,1.20438 3.3116,0.23599 2.52188,-1.37454 l -2.15837,-4.62345 h 4.81656 z" id="path5565" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17453-7);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1.02817345;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
      <ns0:path d="m 736.42336,669.32166 v 16.90341 l 3.8169,-3.72602 2.18109,4.45305 c 0.53423,1.20438 3.3116,0.23599 2.52188,-1.37454 l -2.15837,-4.62345 h 4.81656 z" id="path6242" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17455-1);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1.02817345;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
      <ns0:path d="M 600.56278,703.31514 H 748.51309" id="path9337" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
      <ns0:text id="text9333" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="694.71686" xml:space="preserve"><ns0:tspan id="tspan9335" style="font-size:5.21739101px;line-height:1.25" x="610.1059" y="694.71686" ns2:role="line">Datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:text id="text9341" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="740.54083" y="694.71686" xml:space="preserve"><ns0:tspan id="tspan9343" style="font-size:5.21739101px;line-height:1.25" x="740.54083" y="694.71686" ns2:role="line">1 september 2015, 09:51</ns0:tspan></ns0:text>
      <ns0:text id="text9345" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="717.82251" xml:space="preserve"><ns0:tspan id="tspan9347" style="font-size:5.21739101px;line-height:1.25" x="610.1059" y="717.82251" ns2:role="line">Tidszon</ns0:tspan></ns0:text>
      <ns0:text id="text9349" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="740.54083" y="717.82251" xml:space="preserve"><ns0:tspan id="tspan9351" style="font-size:5.21739101px;line-height:1.25" x="740.54083" y="717.82251" ns2:role="line">CEST (Stockholm, Sverige)</ns0:tspan></ns0:text>
      <ns0:rect height="23.478262" id="rect9353" rx="0" ry="0" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.7453416;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" width="147.9503" x="600.56281" y="742.30591"/>
      <ns0:text id="text9355" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="756.2077" xml:space="preserve"><ns0:tspan id="tspan9357" style="font-size:5.21739101px;line-height:1.25" x="610.1059" y="756.2077" ns2:role="line">Tidsformat</ns0:tspan></ns0:text>
      <ns0:rect height="12.298138" id="rect9363" rx="1.0248625" ry="1.0248625" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.37267077;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" width="38.341366" x="702.89008" y="747.73126"/>
      <ns0:text id="text9359" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="727.87006" y="755.83502" xml:space="preserve"><ns0:tspan id="tspan9361" style="font-size:5.21739101px;line-height:1.25" x="727.87006" y="755.83502" ns2:role="line">24-timmars</ns0:tspan></ns0:text>
      <ns0:path d="m 737.50428,752.6939 -1.96993,1.96993 -1.96993,-1.96993 z" id="rect9365" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" ns2:nodetypes="cccc" ns1:connector-curvature="0"/>
      <ns0:text id="text946" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="541.68079" y="622.67847" xml:space="preserve"><ns0:tspan id="tspan944" style="font-size:5.21739101px;line-height:1.25" x="541.68079" y="622.67847" ns2:role="line">Detaljer</ns0:tspan></ns0:text>
      <ns0:rect height="5.9627328" id="rect948" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.3726708;marker:none;enable-background:new" transform="scale(-1,1)" width="5.9627328" x="-575.56482" y="617.82538"/>
      <ns0:rect height="11.925466" id="rect952" rx="1.4906832" ry="1.4906832" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.3726708;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" width="11.925466" x="566.84741" y="615.02734"/>
      <ns0:g id="g7352" style="display:inline;enable-background:new" transform="matrix(0.37267081,0,0,0.37267081,562.5214,515.34088)" ns1:label="open-menu">
        <ns0:rect height="16" id="rect7354" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" width="16" x="20" y="276"/>
        <ns0:rect height="2.0002136" id="rect7356" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" width="9.9996014" x="23.000198" y="278.99979"/>
        <ns0:rect height="2.0002136" id="rect7358" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" width="9.9996014" x="23.000198" y="282.99979"/>
        <ns0:rect height="2.0002136" id="rect7360" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" width="9.9996014" x="23.000198" y="286.99979"/>
      </ns0:g>
      <ns0:rect height="17.142857" id="rect7822" style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" width="79.006218" x="502.923" y="646.15674"/>
      <ns0:g id="g24827" style="fill:#ffffff;enable-background:new" transform="matrix(0.37267081,0,0,0.37267081,440.68702,454.60394)" ns1:label="preferences-system-time">
        <ns0:circle cx="-9" cy="321" id="path24839" r="7" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#ffffff;stroke-width:2.15384626;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" transform="matrix(0.92857143,0,0,0.92857143,198.85734,238.42857)"/>
        <ns0:path d="m -13.5625,316.46875 3.111031,3.04475 m 0.0029,-0.0135 h 2.948604" id="path25609" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#f7f7f7;stroke-width:1;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" transform="translate(201.0002,217)" ns2:nodetypes="cccc" ns1:connector-curvature="0" ns1:original-d="m -13.5625,316.46875 3.111031,3.04475 m 0.0029,-0.0135 h 2.948604"/>
      </ns0:g>
      <ns0:text id="text7826" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#ffffff;fill-opacity:1;stroke:none" x="536.0907" y="656.21881" xml:space="preserve"><ns0:tspan id="tspan7824" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.21739101px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;fill:#ffffff" x="536.0907" y="656.21881" ns2:role="line">Datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:path d="m 582.12691,611.30064 v 164.9182" id="path7828" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" ns1:connector-curvature="0"/>
      <ns0:rect height="3.3540373" id="rect7830" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" width="17.888199" x="521.92926" y="636.83997"/>
      <ns0:rect height="3.3540373" id="rect7832" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" width="17.888199" x="521.92926" y="670.38031"/>
      <ns0:rect height="3.3540373" id="rect7834" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" width="17.888199" x="521.92926" y="685.28717"/>
      <ns0:rect height="3.3540373" id="rect7836" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" width="28.695652" x="544.28955" y="685.28717"/>
      <ns0:circle cx="511.711" cy="638.71655" id="path7840" r="4.2555118" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle cx="511.711" cy="672.62958" id="circle7842" r="4.2555118" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle cx="511.711" cy="686.79108" id="circle7844" r="4.2555118" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
    </ns0:g>
    <ns0:rect height="29.303314" id="rect3923" rx="14.65165" ry="14.65165" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1" width="53.140442" x="655.56671" y="645.81787"/>
    <ns0:circle cx="693.00433" cy="660.46039" id="path915" r="11.844038" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:16;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
  </ns0:g>
</ns0:svg>
