<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Länka och avlänka kontakter</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="contacts.html" title="Kontakter">Kontakter</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Länka och avlänka kontakter</span></h1></div>
<div class="region">
<div class="contents"></div>
<div id="link-contacts" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Länka kontakter</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan kombinera duplicerade kontakter från din lokala adressbok och nätkonton till en post i <span class="app">Kontakter</span>. Denna funktionen hjälper dig att hålla din adressbok organiserad, med alla detaljer om en kontakt på ett ställe.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Aktivera <span class="em">markeringsläge</span> genom att klicka på bocken ovanför kontaktlistan.</p></li>
<li class="steps"><p class="p">En kryssruta kommer visas bredvid varje kontakt. Kryssa i rutorna vid de kontakter du vill sammanfoga.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Länka</span> för att länka de markerade kontakterna.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="unlink-contacts" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Avlänka kontakter</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan komma att vilja avlänka kontakter om du av misstag länkat samman kontakter som inte ska vara sammanlänkade.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Välj den kontakt du vill avlänka från din kontaktlista.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Redigera</span> i det övre högra hörnet i <span class="app">Contacts</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Länkade kontakter</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Ta bort</span> för att avlänka posten från kontakten.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Stäng</span> när du har avlänkat de poster du vill avlänka.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Färdig</span> för att slutföra redigeringen.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="contacts.html" title="Kontakter">Kontakter</a><span class="desc"> — Kom åt dina kontakter.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
