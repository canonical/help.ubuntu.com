<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Logga ut, stäng av eller växla användare</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Logga ut, stäng av eller växla användare</span></h1></div>
<div class="region">
<div class="contents"><p class="p">När du har använt din dator färdigt kan du stänga av den, försätta din i vänteläge (för att spara ström) eller lämna den på och logga ut.</p></div>
<div id="logout" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Logga ut eller växla användare</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att låta andra användare använda din dator kan du antingen logga ut eller låta dig själv vara inloggad och bara växla användare. Om du växlar användare, kommer alla dina program att fortsätta köra och allting kommer att finnas kvar som där du lämnade det när du logga in igen.</p>
<p class="p">För att <span class="gui">Logga ut</span> eller <span class="gui">Växla användare</span>, klicka på <span class="link"><a href="shell-introduction.html.sv#yourname" title="Du och din dator">systemmenyn</a></span> på höger sida av systemraden, klicka på ditt namn och välj sedan rätt alternativ.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Alternativen <span class="gui">Logga ut</span> och <span class="gui">Växla användare</span> visas bara i meny om du har mer än ett användarkonto på ditt system.</p></div></div></div></div>
</div></div>
</div></div>
<div id="lock-screen" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Lås skärmen</span></h2></div>
<div class="region">
<div class="contents">
<p class="p">Om du ska lämna din dator för en kort stund bör du låsa skärmen för att förhindra andra människor från att nå dina filer eller körande program. När du kommer tillbaka, höj upp gardinen på <span class="link"><a href="shell-lockscreen.html.sv" title="Låsskärmen">låsskärmen</a></span> och mata in ditt lösenord för att logga in igen. Om du inte låser din skärm kommer den automatiskt att låsas efter en viss tid.</p>
<p class="p">För att låsa din skärm, klicka på systemmenyn på höger sida av systemraden och tryck på knappen för att låsa skärmen längst ner på menyn.</p>
<p class="p">När skärmen är låst, kan andra användare logga in på deras egna konton genom att klicka på <span class="gui">Logga in som en annan användare</span> på lösenordsskärmen. Du kan växla tillbaka till ditt skrivbord när de är klara.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="privacy-screen-lock.html.sv" title="Lås automatiskt din skärm">Lås automatiskt din skärm</a><span class="desc"> — Förhindra andra personer från att använda ditt skrivbord när du går iväg från datorn.</span>
</li>
<li class="links ">
<a href="session-screenlocks.html.sv" title="Skärmen låser sig själv allt för snabbt">Skärmen låser sig själv allt för snabbt</a><span class="desc"> — Ändra hur länge det tar innan skärmen låser sig själv i <span class="gui">Sekretessinställningar</span>.</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="suspend" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Vänteläge</span></h2></div>
<div class="region">
<div class="contents">
<p class="p">För att spara ström, försätt din dator i vänteläge när du inte använder den. Om du använder en bärbar dator, kommer GNOME som standard automatiskt att försätta datorn i vänteläge när du stänger locket. Detta sparar tillståndet till din dators minne och stänger av de flesta av datorns funktioner. En väldigt liten del av strömmen används fortfarande i vänteläge.</p>
<p class="p">För att försätta din dator i vänteläge manuellt, klicka på systemmenyn på höger sida av systemraden. Därifrån kan du antingen hålla ner <span class="key"><kbd>Alt</kbd></span>-tangenten och klicka på avstängningsknappen, eller helt enkelt klicka ett långt klick på avstängningsknappen.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="power-batterylife.html.sv" title="Använd mindre ström och förbättra batteridriftstiden">Använd mindre ström och förbättra batteridriftstiden</a><span class="desc"> — Tips på hur du reducerar din dators strömförbrukning.</span>
</li>
<li class="links ">
<a href="power-autosuspend.html.sv" title="Konfigurera automatiskt vänteläge">Konfigurera automatiskt vänteläge</a><span class="desc"> — Konfigurera din dator att automatiskt gå i vänteläge.</span>
</li>
<li class="links ">
<a href="power-suspend.html.sv" title="Vad händer när jag försätter min dator i vänteläge?">Vad händer när jag försätter min dator i vänteläge?</a><span class="desc"> — Vänteläge försätter din dator i ett strömsparläge där den drar mindre ström.</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="shutdown" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Stäng av eller starta om</span></h2></div>
<div class="region">
<div class="contents">
<p class="p">Om du vill stänga av din dator helt eller göra en full omstart, klicka på systemmenyn på höger sida av systemraden och tryck på avstängningsknappen längst ner på menyn. En dialogruta kommer att öppnas som erbjuder dig alternativen att antingen <span class="gui">Starta om</span> eller <span class="gui">Stäng av</span>.</p>
<p class="p">Om det finns andra användare som är inloggade är du kanske inte tillåten att stänga av eller starta om datorn eftersom detta kommer att avsluta deras sessioner. Om du är en administrativ användare kan du bli tillfrågad om ditt lösenord för att stänga av.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan vilja stänga av din dator om du vill flytta den och inte har något batteri, om ditt batteri är lågt eller inte håller laddning bra. En avstängd dator använder också <span class="link"><a href="power-batterylife.html.sv" title="Använd mindre ström och förbättra batteridriftstiden">mindre energi</a></span> än en som är i vänteläge.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="power-batterylife.html.sv" title="Använd mindre ström och förbättra batteridriftstiden">Använd mindre ström och förbättra batteridriftstiden</a><span class="desc"> — Tips på hur du reducerar din dators strömförbrukning.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="shell-overview.html.sv" title="Ditt skrivbord">Ditt skrivbord</a><span class="desc"> — <span class="link"><a href="clock-calendar.html.sv" title="Kalendermöten">Kalender</a></span>, <span class="link"><a href="shell-notifications.html.sv" title="Aviseringar och meddelandefältet">aviseringar</a></span>, <span class="link"><a href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar">tangentbordsgenvägar</a></span>, <span class="link"><a href="shell-windows.html.sv" title="Fönster och arbetsytor">fönster och arbetsytor</a></span>…</span>
</li>
<li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links ">
<a href="power.html.sv" title="Ström och batteri">Ström och batteri</a><span class="desc"> — <span class="link"><a href="power-status.html.sv" title="Kontrollera batteristatus">Batteristatus</a></span>, <span class="link"><a href="power-suspend.html.sv" title="Vad händer när jag försätter min dator i vänteläge?">försätta i vänteläge</a></span>, <span class="link"><a href="power-whydim.html.sv" title="Varför tonas min skärm ner efter ett tag?">skärmtoning</a></span>…</span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="user-autologin.html.sv" title="Logga in automatiskt">Logga in automatiskt</a><span class="desc"> — Ställ in automatisk inloggning när du startar din dator.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p>You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
