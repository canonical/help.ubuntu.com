<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Inledning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="samba.html" title="Samba">Samba</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="samba.html" title="Samba">Föregående</a><a class="nextlinks-next" href="samba-fileserver.html" title="File Server">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Inledning</h1></div>
<div class="region"><div class="contents">
<p class="para">För att använda Ubuntu-system tillsammans med Windowsklienter måste man använda tjänster som är kända i Windowsmiljöer. Sådana tjänster hjälper till att dela data samt information om datorer och användare som är anslutna till nätverket. Dessa tjänster kan delas in tre huvudsakliga kategorier:</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
        <p class="para"><span class="em em-bold emphasis">Fil- och skrivardelning</span>. Använder protokollet Server Message Block (SMB) för att dela filer, mappar, enheter och skrivare i nätverket.</p>
      </li>
<li class="list itemizedlist">
        <p class="para"><span class="em em-bold emphasis">Katalogtjänster</span>. Delar viktig information om datorer och användare i nätverket med hjälp av teknologier som Lightweight Directory Access Protocol (LDAP) och Microsoft <span class="trademark">Active Directory®</span>.</p>
      </li>
<li class="list itemizedlist">
        <p class="para"><span class="em em-bold emphasis">Autentisering och åtkomst</span>. Säkerställer identiteten hos en dator eller användare i ett nätverk och avgör vilken information som dator eller användaren har tillåtelse att nå med hjälp av policys och teknologier som filrättigheter, gruppolicys och autentiseringstjänsten Kerberos.</p>
      </li>
</ul></div>
<p class="para">Dessbättre, kan ditt Ubuntu-system tillhandahålla alla sådana system till Windows-klienter och dela nätverksresurser bland dem. En av de viktigaste programvarorna som ditt Ubuntu-systemet tillhandahåller för Windows-nätverk är Samba-paketet som består av SMB-serverprogram och verktyg.</p>
<p class="para">Detta avsnitt av <span class="phrase">Ubuntu</span> serverguide kommer att introducera några vanliga användningsområden för Samba och hur du installerar och konfigurerar nödvändiga paket. Ytterligare detaljerad dokumentation och information om Samba hittar du på <a href="http://www.samba.org" class="ulink" title="http://www.samba.org">webbplatsen för Samba</a>.</p>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="samba.html" title="Samba">Föregående</a><a class="nextlinks-next" href="samba-fileserver.html" title="File Server">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
