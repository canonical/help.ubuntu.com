<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skicka en fil till en Bluetooth-enhet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="bluetooth.html" title="Bluetooth">Bluetooth</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="sharing.html" title="Sharing">Sharing</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Skicka en fil till en Bluetooth-enhet</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan skicka filer till anslutna Bluetooth-enheter, som mobiltelefoner eller andra datorer. Vissa typer av enheter tillåter inte överföring av filer, eller av vissa filtyper. Du kan skicka filer på tre olika sätt: genom Bluetooth-ikonen i menyraden, från fönstret med Bluetooth-inställningar, eller direkt från filhanteraren.</p>
<p class="p">För att skicka filer direkt från filhanteraren, se <span class="link"><a href="files-share.html" title="Dela ut och överför filer">Dela ut och överför filer</a></span>.</p>
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">Innan du börjar, se till att Bluetooth är aktiverat på din dator. Se zlink xref="bluetooth-turn-on-onff"/&gt;.</p></div></div></div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Skicka filer genom Bluetooth-ikonen</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på Bluetooth-ikonen i menyraden och klicka på <span class="gui">Skicka filer till enhet</span>.</p></li>
<li class="steps">
<p class="p">Välj filen du vill skicka och klicka på <span class="gui">Välj</span>.</p>
<p class="p">För att skicka fler än en fil i en mapp, håll ner <span class="key"><kbd>Ctrl</kbd></span> medan du markerar varje fil.</p>
</li>
<li class="steps">
<p class="p">Markera enheten du vill skicka filerna till och klicka på <span class="gui">Skicka</span>.</p>
<p class="p">Enhetslistan kommer visa både <span class="link"><a href="bluetooth-connect-device.html" title="Anslut din dator till en Bluetooth-enhet">enheter du redan är ansluten till</a></span> och <span class="link"><a href="bluetooth-visibility.html" title="Vad är Bluetooth-synlighet?">synliga enheter</a></span> inom räckhåll. Om du inte redan har anslutit till den markerade enheten kommer du ombes para med enheten när du klickar på <span class="gui">Skicka</span>. Detta kan kräva ytterligare bekräftelse på den andra enheten.</p>
<p class="p">Om det finns många enheter kan du begränsa listan till att bara visa specifika enhetstyper med den utfällbara menyn <span class="gui">Enhetstyper</span>.</p>
</li>
<li class="steps"><p class="p">Ägaren för den mottagande enheten måste oftast trycka på en knapp för att ta emot filen. När ägaren accepterar eller nekar kommer resultat av filöverföringen visas på din skärm.</p></li>
</ol></div>
</div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Skicka filer från Bluetooth-inställningarna</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på Bluetooth-ikonen i menyraden och välj <span class="gui">Bluetooth-inställningar</span>.</p></li>
<li class="steps"><p class="p">Markera enheten du vill skicka filer till från listan till vänster. Listan visar bara enheter du redan har anslutit till. Se <span class="link"><a href="bluetooth-connect-device.html" title="Anslut din dator till en Bluetooth-enhet">Anslut din dator till en Bluetooth-enhet</a></span>.</p></li>
<li class="steps"><p class="p">I enhetsinformationen till höger, klicka <span class="gui">Skicka filer</span>.</p></li>
<li class="steps">
<p class="p">Välj filen du vill skicka och klicka på <span class="gui">Välj</span>.</p>
<p class="p">För att skicka fler än en fil i en mapp, håll ner <span class="key"><kbd>Ctrl</kbd></span> medan du markerar varje fil.</p>
</li>
<li class="steps"><p class="p">Ägaren för den mottagande enheten måste oftast trycka på en knapp för att ta emot filen. När ägaren accepterar eller nekar kommer resultat av filöverföringen visas på din skärm.</p></li>
</ol></div>
</div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="bluetooth.html" title="Bluetooth">Bluetooth</a><span class="desc"> — <span class="link"><a href="bluetooth-connect-device.html" title="Anslut din dator till en Bluetooth-enhet">Anslut</a></span>, <span class="link"><a href="bluetooth-send-file.html" title="Skicka en fil till en Bluetooth-enhet">skicka filer</a></span>, <span class="link"><a href="bluetooth-turn-on-onff.html" title="bluetooth-turn-on-onff">slå på och av</a></span>...</span>
</li>
<li class="links ">
<a href="sharing.html" title="Sharing">Sharing</a><span class="desc"> — 
      <span class="link"><a href="sharing-desktop.html" title="Share your desktop">Desktop sharing</a></span>,
      <span class="link"><a href="files-share.html" title="Dela ut och överför filer">Share files</a></span>…
    </span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-share.html" title="Dela ut och överför filer">Dela ut och överför filer</a><span class="desc"> — För över filer till dina e-postkontakter från filhanteraren.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
