<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ställ in tangentbordsgenvägar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 20.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="keyboard.html.sv" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 20.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="keyboard.html.sv" title="Tangentbord">Tangentbord</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Ställ in tangentbordsgenvägar</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">För att ändra tangenten eller tangenterna som ska tryckas ner för en snabbtangent:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Inställningar</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Inställningar</span>.</p></li>
<li class="steps"><p class="p">Click <span class="gui">Keyboard Shortcuts</span> in the sidebar to open the panel.</p></li>
<li class="steps"><p class="p">Klicka på raden för den önskade åtgärden. Fönstret <span class="gui">Ställ in kortkommando</span> kommer att visas.</p></li>
<li class="steps"><p class="p">Håll ner den önskade tangentkombinationen eller tryck på <span class="key"><kbd>Backsteg</kbd></span> för att återställa, eller tryck på <span class="key"><kbd>Esc</kbd></span> för att avbryta.</p></li>
</ol></div></div></div>
</div>
<section id="defined"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Fördefinierade tangentbordsgenvägar</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Det finns ett antal förkonfigurerade snabbtangenter som kan ändras, grupperade i dessa kategorier:</p>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">Programstartare</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Hem-mapp</p></td>
<td><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-folder.svg" class="media media-inline" alt="Explorer key symbol"></span></span> eller <span class="media"><span class="media media-image"><img src="figures/keyboard-key-computer.svg" class="media media-inline" alt="Explorer key symbol"></span></span> eller <span class="key"><kbd>Utforskare</kbd></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Starta kalkylator</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-calculator.svg" class="media media-inline" alt="Calculator key symbol"></span></span> eller <span class="key"><kbd>Kalkylator</kbd></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Starta e-postklient</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-mail.svg" class="media media-inline" alt="Mail key symbol"></span></span> eller <span class="key"><kbd>E-post</kbd></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Start hjälpläsare</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Starta webbläsare</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-world.svg" class="media media-inline" alt="WWW key symbol"></span></span> eller <span class="media"><span class="media media-image"><img src="figures/keyboard-key-home.svg" class="media media-inline" alt="WWW key symbol"></span></span> eller <span class="key"><kbd>WWW</kbd></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Sök</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-search.svg" class="media media-inline" alt="Search key symbol"></span></span> eller <span class="key"><kbd>Sök</kbd></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Inställningar</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Verktyg</kbd></span></p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">Navigering</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Göm alla normala fönster</p></td>
<td><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta en arbetsyta uppåt</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Up</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta en arbetsyta nedåt</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Down</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster en skärm nedåt</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span>+<span class="key"><kbd>↓</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster en skärm åt vänster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>←</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster en skärm åt höger</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>→</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster en skärm uppåt</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>↑</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster en arbetsyta nedåt</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Down</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster en arbetsyta uppåt</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Up</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster till sista arbetsyta</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>End</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster till arbetsyta 1</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Home</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster till arbetsyta 2</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster till arbetsyta 3</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster till arbetsyta 4</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla program</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla systemkontroller</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla systemkontroller omedelbart</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Esc</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla till sista arbetsyta</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>End</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla till arbetsyta 1</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Home</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla till arbetsyta 2</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla till arbetsyta 3</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla till arbetsyta 4</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla mellan fönster</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla fönster omedelbart</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Esc</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla direkt mellan fönster i ett program</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F6</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla mellan fönster i ett program</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">Skärmbilder</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Kopiera en skärmbild av ett fönster till urklipp</p></td>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Kopiera en skärmbild av ett område till urklipp</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Kopiera en skärmbild till urklipp</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Spela in en kort skärminspelning</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>R</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Spara en skärmbild av ett fönster till Bilder</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Spara en skärmbild av ett område till Bilder</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Spara en skärmbild till Bilder</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Print</kbd></span></p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">Ljud och media</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Mata ut</p></td>
<td><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-eject.svg" class="media media-inline" alt="Eject key symbol"></span></span> (Mata ut)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Starta mediaspelare</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-media.svg" class="media media-inline" alt="Media key symbol"></span></span> (Ljud media)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Nästa spår</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-next.svg" class="media media-inline" alt="Next key symbol"></span></span> (Ljud nästa)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Pausa uppspelning</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-pause.svg" class="media media-inline" alt="Pause key symbol"></span></span> (Ljud pausa)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Spela (eller spela/pausa)</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-play.svg" class="media media-inline" alt="Play key symbol"></span></span> (Ljud spela upp)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Föregående spår</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-previous.svg" class="media media-inline" alt="Previous key symbol"></span></span> (Ljud föregående)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Stoppa uppspelning</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-stop.svg" class="media media-inline" alt="Stop key symbol"></span></span> (Ljud stoppa)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Sänk volymen</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-voldown.svg" class="media media-inline" alt="Volume Down key symbol"></span></span> (Ljud sänk volym)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Tyst</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-mute.svg" class="media media-inline" alt="Mute key symbol"></span></span> (Ljud stäng av)</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Höj volymen</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/keyboard-key-volup.svg" class="media media-inline" alt="Volume Up key symbol"></span></span> (Ljud höj volym)</p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">System</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Skifta fokus till den aktiva aviseringen</p></td>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>N</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Låsskärmen</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>L</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Logga ut</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Delete</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Öppna programmenyn</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>F10</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Återställ tangentbordsgenvägarna</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Esc</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Visa alla program</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>A</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Visa aktivitetsöversiktsvyn</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F1</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Visa aviseringslistan</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>V</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Visa översiktsvyn</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>S</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Visa rutan kör ett kommando</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F2</kbd></span></span></p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">Skriva</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Byt till nästa inmatningskälla</p></td>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">By till föregående inmatningskälla</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span></p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">Hjälpmedel</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Minska textstorleken</p></td>
<td><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Hög kontrast på eller av</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Öka textstorleken</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Aktivera eller inaktivera skärmtangentbord</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Aktivera eller inaktivera skärmläsare</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>S</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Aktivera eller inaktivera zoom</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>8</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Zooma in</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>=</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Zooma ut</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>-</kbd></span></span></p></td>
</tr>
</table></div>
</div>
</div>
<div class="table ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-table"><h3><span class="title">Fönster</span></h3></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p">Aktivera fönstermenyn</p></td>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Stänga fönster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F4</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Göm fönster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>H</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Sänk fönstret under andra fönster</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Maximera fönster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>↑</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Maximera fönster horisontellt</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Maximera fönster vertikalt</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Flytta fönster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F7</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Höj fönstret över andra fönster</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Höj fönstret om det skyms, sänk det annars</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Storleksändra fönster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F8</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Återställ fönster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>↓</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla helskärmsläge</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla maximeringstillstånd</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F10</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Växla fönster på alla arbetsytor eller bara en</p></td>
<td style="border-top-style: solid;"><p class="p">Inaktiverad</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Vy delad till vänster</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>←</kbd></span></span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Vy delad till höger</p></td>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>→</kbd></span></span></p></td>
</tr>
</table></div>
</div>
</div>
</div></div>
</div></section><section id="custom"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Anpassade genvägar</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">För att skapa dina egna snabbtangenter för program i inställningarna för <span class="app">Tangentbord</span>:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på knappen <span class="gui">+</span>. Fönstret <span class="gui">Lägg till anpassat kortkommando</span> kommer att visas.</p></li>
<li class="steps"><p class="p">Mata in ett <span class="gui">Namn</span> för att identifiera genvägen och ett <span class="gui">Kommando</span> för att köra ett program. Om du till exempel ville att genvägen ska öppna <span class="app">Rhythmbox</span>, kan du namnge den <span class="input">Musik</span> och använda kommandot <span class="input">rhythmbox</span>.</p></li>
<li class="steps"><p class="p">Klicka på raden som just lades till. Då fönstret <span class="gui">Ställ in anpassat kortkommando</span> öppnas, tryck ner den önskade tangentkombinationen för kortkommandot.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Lägg till…</span>.</p></li>
</ol></div></div></div>
<p class="p">Kommandonamnet som du matade in bör vara ett giltigt systemkommando. Du kan kontrollera att kommandot fungerar genom att öppna en Terminal och skriva in det där. Kommandot som öppnar ett program kan inte ha samma namn som programmet själv.</p>
<p class="p">Om du vill ändra kommandot som är associerat med en anpassad tangentbordsgenväg, dubbelklicka på genvägens <span class="em">namn</span>. Fönstret <span class="gui">Ställ in anpassat kortkommando</span> kommer att visas och du kan redigera kommandot.</p>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="keyboard.html.sv" title="Tangentbord">Tangentbord</a><span class="desc"> — <span class="link"><a href="keyboard-layouts.html.sv" title="Använd alternativa tangentbordslayouter">Tangentbordslayouter</a></span>, <span class="link"><a href="keyboard-cursor-blink.html.sv" title="Få tangentbordsmarkören att blinka">markörblinkning</a></span>, <span class="link"><a href="a11y.html.sv#mobility" title="Rörelsehinder">tangentbordshjälpmedel</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar">Användbara tangentbordsgenvägar</a><span class="desc"> — Ta sig runt på skrivbordet med hjälp av tangentbordet.</span>
</li></ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
