<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ditt skrivbord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Ditt skrivbord</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-introduction.html.sv" title="Introduktion till GNOME"><span class="title">Introduktion till GNOME</span><span class="linkdiv-dash"> — </span><span class="desc">En visuell introduktion till ditt skrivbord, systemraden, och översiktsvyn <span class="gui">Aktiviteter</span>.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-exit.html.sv" title="Logga ut, stäng av eller växla användare"><span class="title">Logga ut, stäng av eller växla användare</span><span class="linkdiv-dash"> — </span><span class="desc">Lär dig hur du lämnar ditt användarkonto genom att logga ut, växla användare, och så vidare.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="shell-apps-open.html.sv" title="Starta program"><span class="title">Starta program</span><span class="linkdiv-dash"> — </span><span class="desc">Starta program från översiktsvyn <span class="gui">Aktiviteter</span>.</span></a></div></div>
</div></div></div></div>
<div id="desktop" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Anpassa ditt skrivbord</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-notifications.html.sv" title="Aviseringar och meddelandefältet"><span class="title">Aviseringar och meddelandefältet</span><span class="linkdiv-dash"> — </span><span class="desc">Meddelanden visas längst upp på skärmen för att berätta för dig när vissa händelser inträffar.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="clock-calendar.html.sv" title="Kalendermöten"><span class="title">Kalendermöten</span><span class="linkdiv-dash"> — </span><span class="desc">Visa dina möten i kalenderområdet i toppen på skärmen.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="shell-apps-favorites.html.sv" title="Nåla fast dina favoritprogram i snabbstartspanelen"><span class="title">Nåla fast dina favoritprogram i snabbstartspanelen</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till (eller ta bort) ofta använda programikoner från snabbstartspanelen.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="apps" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Program och fönster</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar"><span class="title">Användbara tangentbordsgenvägar</span><span class="linkdiv-dash"> — </span><span class="desc">Ta sig runt på skrivbordet med hjälp av tangentbordet.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-windows.html.sv" title="Fönster och arbetsytor"><span class="title">Fönster och arbetsytor</span><span class="linkdiv-dash"> — </span><span class="desc">Flytta och organisera dina fönster.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-lockscreen.html.sv" title="Låsskärmen"><span class="title">Låsskärmen</span><span class="linkdiv-dash"> — </span><span class="desc">Den dekorativa och funktionella låsskärmen förmedlar användbar information.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="startup-applications.html.sv" title="Uppstartsprogram"><span class="title">Uppstartsprogram</span><span class="linkdiv-dash"> — </span><span class="desc">Välj vilka program som skall startas när du loggar in.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="status-icons.html.sv" title="Vad betyder ikonerna i systemraden?"><span class="title">Vad betyder ikonerna i systemraden?</span><span class="linkdiv-dash"> — </span><span class="desc">Förklarar innebörden av ikonerna som finns i den högra delen av systemraden.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-windows-switching.html.sv" title="Växla mellan fönster"><span class="title">Växla mellan fönster</span><span class="linkdiv-dash"> — </span><span class="desc">Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span>.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
