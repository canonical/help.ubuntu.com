<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Hjälpmedel</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 25.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Hjälpmedel</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Systemet inkluderar hjälpmedelsteknik för att stödja användare med olika typer av funktionshinder och speciella behov och för att interagera med vanliga hjälpmedelsenheter. En hjälpmedelsmeny kan läggas till i systemraden och lätt ge tillgång till många av hjälpmedelsfunktionerna.</p>
<div class="links topiclinks"><div class="inner"><div class="region"><div class="links-divs"><div class="linkdiv "><a class="linkdiv" href="a11y-icon.html.sv" title="Hitta hjälpmedelsmenyn"><span class="title">Hitta hjälpmedelsmenyn</span><span class="linkdiv-dash"> — </span><span class="desc">Hjälpmedelsmenyn är ikonen i systemraden som ser ut som en person.</span></a></div></div></div></div></div>
</div>
<section id="vision"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Synnedsättningar</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h3><span class="title">Blindhet</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="a11y-screen-reader.html.sv" title="Högläsning av skärmen">Högläsning av skärmen</a><span class="desc"> — Använd skärmläsaren <span class="app">Orca</span> för att läsa upp användargränssnittet.</span>
</li>
<li class="links ">
<a href="a11y-braille.html.sv" title="Läs skärmen med punktskrift">Läs skärmen med punktskrift</a><span class="desc"> — Använd skärmläsaren <span class="app">Orca</span> med en uppdateringsbar punktskriftsskärm.</span>
</li>
</ul></div>
</div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h3><span class="title">Nedsatt syn</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="keyboard-cursor-blink.html.sv" title="Få tangentbordsmarkören att blinka">Få tangentbordsmarkören att blinka</a><span class="desc"> — Få insättningspunkten att blinka och kontrollera hur snabbt den blinkar.</span>
</li>
<li class="links ">
<a href="a11y-mag.html.sv" title="Förstora en del av skärmen">Förstora en del av skärmen</a><span class="desc"> — Zooma in på din skärm så att det är enklare att se saker.</span>
</li>
<li class="links ">
<a href="a11y-contrast.html.sv" title="Justera kontrasten">Justera kontrasten</a><span class="desc"> — Gör fönster och knappar på skärmen mer (eller mindre) tydliga så de är enklare att se.</span>
</li>
<li class="links ">
<a href="a11y-font-size.html.sv" title="Ändra textstorlek på skärmen">Ändra textstorlek på skärmen</a><span class="desc"> — Använd större typsnitt för att göra text enklare att läsa.</span>
</li>
</ul></div>
</div></div>
</div></div>
</div></section><section id="sound"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Hörselnedsättningar</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><ul><li class="links ">
<a href="a11y-visualalert.html.sv" title="Blinka skärmen vid larmljud">Blinka skärmen vid larmljud</a><span class="desc"> — Aktivera visuella larm för att få skärmen eller fönstret att blinka när ett larmljud spelas.</span>
</li></ul></div></div></div></div></div>
</div></section><section id="mobility"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Rörelsehinder</span></h2></div>
<div class="region">
<div class="contents pagewide">
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h3><span class="title">Musförflyttning</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="mouse-sensitivity.html.sv" title="Justera hastigheten för musen och styrplattan">Justera hastigheten för musen och styrplattan</a><span class="desc"> — Ändra hur snabbt markören flyttar sig när du använder din mus eller styrplatta.</span>
</li>
<li class="links ">
<a href="mouse-mousekeys.html.sv" title="Klicka och flytta muspekaren med det numeriska tangentbordet">Klicka och flytta muspekaren med det numeriska tangentbordet</a><span class="desc"> — Aktivera mustangenter för att styra musen med det numeriska tangentbordet.</span>
</li>
</ul></div>
</div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h3><span class="title">Klicka och dra</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="mouse-doubleclick.html.sv" title="Justera hastigheten för dubbelklick">Justera hastigheten för dubbelklick</a><span class="desc"> — Styr hur snabbt du behöver trycka på musknappen en andra gång för att dubbelklicka.</span>
</li>
<li class="links ">
<a href="a11y-right-click.html.sv" title="Simulera ett högerklick">Simulera ett högerklick</a><span class="desc"> — Tryck och håll kvar vänstra musknappen för att högerklicka.</span>
</li>
<li class="links ">
<a href="a11y-dwellclick.html.sv" title="Simulera klick genom att sväva ovanför">Simulera klick genom att sväva ovanför</a><span class="desc"> — Funktionen <span class="gui">Uppehållsklick</span> (svävningsklick) låter dig klicka genom att hålla muspekaren stilla.</span>
</li>
</ul></div>
</div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h3><span class="title">Användning av tangentbord</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="a11y-stickykeys.html.sv" title="Aktivera klistriga tangenter">Aktivera klistriga tangenter</a><span class="desc"> — Mata in snabbtangenter en tangent i taget i stället för att hålla ner alla tangenterna på en gång.</span>
</li>
<li class="links ">
<a href="a11y-bouncekeys.html.sv" title="Aktivera tangentstuds">Aktivera tangentstuds</a><span class="desc"> — Ignorera snabbt upprepade tangenttryckningar på samma tangent.</span>
</li>
<li class="links ">
<a href="a11y-slowkeys.html.sv" title="Aktivera tröga tangenter">Aktivera tröga tangenter</a><span class="desc"> — Aktivera en fördröjning mellan tangenttryckning till det att bokstaven syns på skärmen.</span>
</li>
<li class="links ">
<a href="keyboard-osk.html.sv" title="Använd ett skärmtangentbord">Använd ett skärmtangentbord</a><span class="desc"> — Använd ett skärmtangentbord för att mata in text genom att klicka på knappar med musen eller en pekskärm.</span>
</li>
<li class="links ">
<a href="keyboard-repeat-keys.html.sv" title="Hantera upprepade tangenttryckningar">Hantera upprepade tangenttryckningar</a><span class="desc"> — Få tangentbordet att inte upprepa bokstäver när du håller ner en tangent, eller ändra fördröjningen och hastigheten på upprepande tangenter.</span>
</li>
<li class="links ">
<a href="keyboard-nav.html.sv" title="Tangentbordsnavigation">Tangentbordsnavigation</a><span class="desc"> — Använd program och skrivbordet utan en mus.</span>
</li>
</ul></div>
</div></div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="keyboard-key-menu.html.sv" title="Vad är Windows-tangenten?">Vad är <span class="key"><kbd>Windows</kbd></span>-tangenten?</a><span class="desc"> — Tangenten <span class="key"><kbd>Meny</kbd></span> startar en snabbvalsmeny med tangentbordet snarare än med ett högerklick.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
