<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använd Synaptic för en mer avancerad programhantering</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="addremove.html.sv" title="Installera &amp; ta bort mjukvara">Lägg till/ta bort program</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Använd Synaptic för en mer avancerad programhantering</span></h1></div>
<div class="region">
<div class="contents">
<p class="p"><span class="app">Synaptic pakethanterare</span> är kraftfullare och kan hantera en del programhanteringsuppgifter som <span class="app">Programvara för Ubuntu</span> inte kan. Synaptics gränssnitt är mera komplicerat och stödjer inte nyare funktioner i <span class="app">Programvara för Ubuntu</span> såsom betygssättning och kommentarer, och rekommenderas därför inte för nya Ubuntu-användare.</p>
<p class="p">Synaptic är inte installerat som standard, men du kan <span class="link"><a href="https://apps.ubuntu.com/cat/applications/synaptic" title="https://apps.ubuntu.com/cat/applications/synaptic">installera</a></span> det från Ubuntus paketförråd.</p>
</div>
<div id="install-software-with-synaptic" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Installera program med Synaptic</span></h2></div>
<div class="region"><div class="contents">
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna <span class="app">Synaptic</span> via sökraden för <span class="em">Aktiviteter</span>. Du behöver ange ditt lösenord i fönstret <span class="gui">Autentisera</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Sök</span> för att söka efter ett program, eller klicka på <span class="gui">Sektioner</span> och gå igenom de olika kategorierna.</p></li>
<li class="steps"><p class="p">Högerklicka på programmet du vill installera och välj <span class="gui">Markera för installation</span>.</p></li>
<li class="steps"><p class="p">Om du ombes markera ytterligare ändringar, klicka på <span class="gui">Markera</span>.</p></li>
<li class="steps"><p class="p">Markera något annat program som du vill installera.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Tillämpa</span>, och klicka sedan på <span class="gui">Tillämpa</span> i fönstret som visas. Programmen du valde kommer laddas ner och installeras.</p></li>
</ol></div></div></div>
<p class="p">För mer information om hur du använder <span class="app">Synaptic</span> hänvisar vi till <span class="link"><a href="https://help.ubuntu.com/community/SynapticHowto" title="https://help.ubuntu.com/community/SynapticHowto">Synaptics handledning</a></span>.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="addremove.html.sv" title="Installera &amp; ta bort mjukvara">Installera &amp; ta bort mjukvara</a><span class="desc"> — <span class="link"><a href="addremove-install.html.sv" title="Installera fler program">Installera program</a></span>, <span class="link"><a href="addremove-remove.html.sv" title="Ta bort ett program">ta bort program</a></span>, <span class="link"><a href="addremove-sources.html.sv" title="Lägg till fler programförråd">lägg till förråd</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="addremove-install.html.sv" title="Installera fler program">Installera fler program</a><span class="desc"> — Använd <span class="app">Programvara för Ubuntu</span> för att lägga till program och göra Ubuntu mer användbart.</span>
</li>
<li class="links ">
<a href="addremove-remove.html.sv" title="Ta bort ett program">Ta bort ett program</a><span class="desc"> — Ta bort program som du inte längre använder.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
