<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Varför känns inte min musikspelare igen när jag ansluter den?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Varför känns inte min musikspelare igen när jag ansluter den?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om din musikspelare (MP3-spelare mm.) ansluts till datorn men inte visas i ditt musikprogram kan den ha felaktigt identifierats som något annat än en musikspelare.</p>
<p class="p">Testa att koppla bort spelaren och sedan ansluta den igen. Om det inte hjälper, <span class="link"><a href="files-browse.html" title="Bläddra bland filer och mappar">öppna filhanteraren</a></span>. Du bör se spelaren i listan under <span class="gui">Enheter</span> i sidoraden - klicka på den för att öppna mappen för musikspelaren. Klicka nu på <span class="guiseq"><span class="gui">Fil</span> ▸ <span class="gui">Nytt dokument</span> ▸ <span class="gui">Tomt dokument</span></span>, skriv <span class="input">.is_audio_player</span> och tryck <span class="key"><kbd>Retur</kbd></span> (punkten och understrecken är viktiga, och allt ska skrivas med små bokstäver). Filen upplyser din dator om att enheten är en musikspelare.</p>
<p class="p">Leta nu efter musikspelaren i filhanterarens sidorad och mata ut den (högerklicka och klicka på <span class="gui">Mata ut</span>). Koppla ur den, och anslut den sedan på nytt. Den här gången bör den identifieras som en musikspelare av ditt musikprogram. Om inte, testa att stänga musikprogrammet och starta det på nytt.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Dessa instruktioner kommer inte fungera för iPod och vissa andra musikspelare. De bör fungera om din spelare är en <span class="em">USB-masslagringsenhet</span>; det bör stå i användarhandboken om spelaren är en sådan.</p></div></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">När du tittar i musikspelarens mapp igen, ser du inte filen <span class="input">.is_audio_player</span>. Detta beror på att punkten i filnamnet talar om för filhanteraren att filen ska döljas. Du kan kontrollera att den fortfarande finns genom att klicka på <span class="guiseq"><span class="gui">Visa</span> ▸ <span class="gui">Visa dolda filer</span></span>.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="music-player-newipod.html" title="Min nya iPod fungerar inte">Min nya iPod fungerar inte</a><span class="desc"> — Helt nya iPods måste ställas in via iTunes-programvaran innan du kan använda dem.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
