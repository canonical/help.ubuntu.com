<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skriv filer till en cd- eller dvd-skiva</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Skriv filer till en cd- eller dvd-skiva</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan spara filer på en blank skiva genom att använda <span class="gui">Cd/dvd-skaparen</span>. Alternativet att skapa en cd eller dvd kommer att synas i filhanteraren så snart du placerat en cd i din cd/dvd-skrivare. Filhanteraren låter dig överföra filer till andra datorer eller utföra <span class="link"><a href="backup-why.html" title="Säkerhetskopiera dina viktiga filer">säkerhetskopiering</a></span> genom att spara filer på en blank skiva. För att skriva filer till en cd eller dvd:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Mata in en tom skiva i din cd-/dvd-brännarenhet.</p></li>
<li class="steps">
<p class="p">I aviseringen <span class="gui">Tom cd/dvd-r-skiva</span> soom visas i botten på skärmen, välj <span class="gui">Öppna med Cd/dvd-skaparen</span>. Mappfönstret <span class="gui">Cd/dvd-skaparen</span> kommer att öppnas.</p>
<p class="p">(Du kan också klicka på <span class="gui">Tom cd/dvd-r skiva</span> under <span class="gui">Enheter</span> i filhanterarens sidopanel.)</p>
</li>
<li class="steps"><p class="p">I fältet <span class="gui">Skivnamn</span>, skriv in ett namn på skivan.</p></li>
<li class="steps"><p class="p">Dra eller kopiera de önskade filerna in i fönstret.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Skriv till skiva</span>.</p></li>
<li class="steps">
<p class="p">Under <span class="gui">Välj en skiva att skriva till</span>, välj den tomma skivan.</p>
<p class="p">(Du kan välja <span class="gui">Avbildningsfil</span> istället. Detta kommer att spara filerna i en <span class="em">skivavbildning</span> vilken kommer att sparas på din dator. Du kan sedan bränna den skivavbildningen på en tom skiva vid ett senare tillfälle.)</p>
</li>
<li class="steps"><p class="p">Klicka på <span class="gui">Egenskaper</span> om du vill justera brännhastighet, plats för tillfälliga filer eller andra inställningar. Standardinställningarna bör duga fint.</p></li>
<li class="steps">
<p class="p">Klicka på knappen <span class="gui">Bränn</span> för att börja skrivningen.</p>
<p class="p">Om <span class="gui">Bränn flera kopior</span> markeras kommer du tillfrågas om ytterligare skivor.</p>
</li>
<li class="steps"><p class="p">När skivbränningen är färdig kommer skivan matas ut automatiskt. Välj <span class="gui">Gör fler kopior</span> eller <span class="gui">Stäng</span> för att avsluta.</p></li>
</ol></div></div></div>
</div>
<div id="problem" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Om skivan inte brändes korrekt</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Ibland bränns skivan inte korrekt, och du kommer inte kunna se filerna på skivan när du matar in den i en dator.</p>
<p class="p">Om detta händer, försöka att bränna skivan igen men använd en lägre brännhastighet, till exempel 12x istället för 48x. Att bränna på lägre hastigheter är mer tillförlitligt. Du kan välja hastighet genom att klicka på <span class="gui">Egenskaper</span> i fönstret <span class="gui">Cd/dvd-skaparen</span>.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
