<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Behöver jag ett anti-virusprogram?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-security.html" title="Trygghet på internet">Trygghet på internet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Behöver jag ett anti-virusprogram?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du är van vid Windows eller Mac OS är du förmodligen också van vid att konstant ha ett aktivt körande anti-virusprogram hela tiden. Anti-virusprogram kör i bakgrunden, och letar konstant efter datorvirus som kan leta sig in i din dator och orsaka problem.</p>
<p class="p">Anti-virusprogram finns för Linux, men du behöver troligtvis inte använda dem. Virus som påverkar Linux är fortfarande mycket sällsynta. Vissa menar att det här beror på att Linux inte används i lika stor utsträckning som de andra operativsystemen, så ingen bryr sig om att skriva virus för det. Andra hävdar att Linux är mer säkert till sin natur, och säkerhetsproblem som virus kan använda sig av lagas mycket snabbt.</p>
<p class="p">Vad sanningen än är, så är Linux-virus så sällsynta att du nog inte behöver oroa dig i dagsläget.</p>
<p class="p">Om du vill vara ännu mer säker, eller om du vill leta efter virus i filer som du skickar mellan dig själv och personer som använder Windows eller Mac OS, kan du så klart installera anti-virusprogram. Sök i <span class="app">Programvara för Ubuntu</span> där ett antal program finns tillgängliga.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-security.html" title="Trygghet på internet">Trygghet på internet</a><span class="desc"> — <span class="link"><a href="net-antivirus.html" title="Behöver jag ett anti-virusprogram?">Antivirusprogram</a></span>, <span class="link"><a href="net-firewall-on-off.html" title="Kontrollera nätverkstrafiken till och från din dator">grundläggande brandväggar</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-email-virus.html" title="Behöver jag söka igenom min e-post efter virus?">Behöver jag söka igenom min e-post efter virus?</a><span class="desc"> — Virus kommer sannolikt inte infektera din dator, men kan infektera datorerna hos personer du skickar e-post till.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
