<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Lås automatiskt din skärm</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="prefs-display.html" title="Visning och skärm">Visning och skärm</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Lås automatiskt din skärm</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">När du går ifrån din dator bör du <span class="link"><a href="shell-exit.html#lock-screen" title="Lås skärmen">låsa skärmen</a></span> för att hindra andra från att använda ditt skrivbord och komma åt dina filer. Du kommer fortfarande vara inloggad, och alla dina program kommer fortfarande köras, men du måste skriva in ditt lösenord igen innan du kan fortsätta använda datorn. Du kan låsa skärmen manuellt, men du kan också låta skärmen låsas automatiskt.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="em">Systemmenyn</span> <span class="media"><span class="media media-image"><img src="figures/system-devices-panel.svg" class="media media-inline" alt="Kugghjulsikon"></span></span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Ljusstyrka &amp; skärmlås</span>.</p></li>
<li class="steps"><p class="p">Se till att <span class="gui">Lås</span> är aktiverat, och välj sedan en tidsgräns från den utfällbara listan nedanför. Skärmen kommer automatiskt låsas efter att du varit inaktiv såpass länge. Du kan också välja <span class="gui">Skärmen stängs av</span> för att låsa skärmen efter att den automatiskt stängs av, vilket styrs av den utfällbara listan <span class="gui">Stäng av skärmen när inaktiv i</span> ovanför.</p></li>
</ol></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs-display.html" title="Visning och skärm">Visning och skärm</a><span class="desc"> — <span class="link"><a href="look-background.html" title="Byt skrivbordsbakgrund">Bakgrund</a></span>, <span class="link"><a href="look-resolution.html" title="Ändra storlek och rotation för skärmen">storlek och orientering</a></span>, <span class="link"><a href="display-dimscreen.html" title="Ställ in skärmens ljusstyrka">ljusstyrka</a></span>...</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="shell-exit.html#lock-screen" title="Lås skärmen">Lås skärmen</a></li>
<li class="links ">
<a href="session-screenlocks.html" title="Skärmen låser sig själv allt för snabbt">Skärmen låser sig själv allt för snabbt</a><span class="desc"> — Ändra hur lång tid det får gå innan skärmen låses i inställningarna för <span class="gui">Ljusstyrka &amp; Lås</span>.</span>
</li>
<li class="links ">
<a href="display-dimscreen.html" title="Ställ in skärmens ljusstyrka">Ställ in skärmens ljusstyrka</a><span class="desc"> — Minska skärmens ljusstyrka för att spara energi, eller öka ljusstyrkan för att göra den mer lättläst i starkt ljus.</span>
</li>
<li class="links ">
<a href="security-settings.html" title="Säkerhet &amp; sekretess">Säkerhet &amp; sekretess</a><span class="desc"> — Ändra några säkerhets- och sekretessinställningar.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
