�PNG

   IHDR  v      ә   �zTXtRaw profile type exif  x�mP�� ���/�iR�t�p���!s������&-�W�jj�t\�Ʉ:y�U�T/:P�K�8��aO�N=/�+yD�è�3�]��߿��!q{Y	����oa��>��xE_m�:+�߽���^�a>�ĂIt c
�G ���%��.*5+�����	xY�Y��0U  �iCCPICC profile  x�}�=H�@�_S�"�q�P����U(B�P+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�F�iV�,�鶙N&�lnU�"�D0Qf�1'I)���{�z�Y���}j�b@@$�e�ioOo��}�(+�*�9�I$~�����ό���<q�X,v����dj�S�1U�)_�z�r��Uj�uO��p^_Y�:�a$��%H���2*��U'�B��>�!�/�K!W��B������w�Var�K
'����B�@��8�ǎ�<������W��'���;����붦��;���!��+i
��~Fߔ"�@��[k�@��J� ��h���}����ۿgZ�� ��r�(˞�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:c5a0a3f4-0793-4bfe-aabf-9c692020ffdc"
   xmpMM:InstanceID="xmp.iid:f6c97e1f-7707-48b7-bf96-d4bc8a0bd00f"
   xmpMM:OriginalDocumentID="xmp.did:1af17f3a-e109-47af-8ea9-43c3ba983090"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679601346795058"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T20:55:46+01:00"
   xmp:ModifyDate="2023:03:23T20:55:46+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:6e1a15d6-7c40-41df-8c06-9a485e1409dd"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T20:55:46+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>�z
�   	pHYs  �  ��+   tIME�8zw   tEXtComment Created with GIMPW�  �IDATx���{TW~�;3z���$� �H�;`����m��c��c��89�I�M�i��{�M�I����n��m���O�d��['��X�� #!�'BB��cn�Pc���������j�8�;�#      �c�      �	C      ���     s1DL     0�     ����ϟ;O�h��^�_VQ������/]�\UY)
g1�B9    ����ׯ���d2�*++�(/�}ݯ;�&Ij�E��d2II~˝9�p(4r�\{������FOOK����1����X,�AH���������><|��+�L�	ӊ�H$���v����,G    ��@ p��+
����z=I�~����w,�ŋ-b��s�b(2������*Uaa!EQ!��e�q��f/)+�r��UI$��������D"q���!���fb�hn��H$R�!D���W����=�v=����D��������"� f��������[m�=�l8v�\o��+����g��uӨ��546:#2����K��~��p���.\�xQ���9sv���!���̙�ŋo�!����&�-���+    �7�O>�,
���'���T"���ys����g�F������m����GG��D���E*�*�r������x���n��V\��L���;7�(6��r��~��	.��y�t����K�vLF#�.\���!���j���Բ�lo���Mo��ꌌ����!�ȈT*�)����>���+O�zB$557o{x[�<�DS3���p�l�B���$I��5�kKK��w_(
���d��q��J�\��z�lvaQ!�ǋ���e<4.
eR)����A�@�R)�`�(3/7���Y��X|tt�/�+
��=����YeA�su9�֭��b��~������b�1f�^���P<�h�*�����;.��l�$��b��#2�,//�apoo�X`L�P�՚X����1�P~~��	   �� ЎG��rL,3���
+++*++BK�J߭�[����b!����6L�Q���rt�`������Z�6����A�X�����oR,��t��z�Xtk�[�<�j���tvv.4���

�7oڔL2����-YZ��p����v�D�`p���U�V!��j�3��A.���={�x�{s�����拕�k~���>���Or���6�r������0�0M�m��@����p8�w�NwǺ���_}��c;7nX��m�����8�~����?y�TUU�y3��;���c�1fs8\c|�ܹ+W�B�бc�*��������m�nmk3�L*���ŋk׬V)U|���`Xh4fffv^31s���7,��8}�K�۝��o2�A^^��f��u�S�����9�5� ���0�a��hpp���?::z����^x!��hz|<��O��b��TJe$��͹z����Zm[[���7sy�_��VQQ��Ź��s�%    �w��*1����L-2�mm�����
N��ݺ���R�������r�'��v=�P(4�L�D���-n.)Y���<�r���(
�(�-�ѨP(���v����cL��J�t9]kW�����?������D!<�0��h���9'��Խ���뽵���-]]]S%;w��h��+vuwޒD�L&3���O��MQT4���.����UWWc�5�O_�IV�c\]]u��!�χ�~ƈ9�����j�v�t��'_�'�e%%�7o"I�DS�R�ܼiS�����%}�ӧO���?�H$$I&I�p�N���m|� !�a���X�a����e�����U+�JE{�����v���߭��w��v�L&����z�~xx8u�a45M ��o?�9ts�����9��:����Y���t�,����>���֭]�P��nwWWWYY�\.ߺe�L&���   ����r�Y,k֬I-vtt��G�x�-�d25]!,��7n܀1~��n\�A,y<�����+W�_�nl,@�t����d1Bh���55�'�����^3�v�z�a�t��p8�r��O�tzzzYY)��d2�\��{����֜����ۗ.YB�Ĝ���Ȉ��u��]�`Bh�р�Z�#N���XQa�L�21�ܖ I��(*�L��r�%3�1�ڀ���e�*&?�d0�0�]:|����X�V��4ui�:6��0���E%�������#IB��K$��3�HH$R�$�lFc���X,6A �o��Ͽ��~�� �EQAȤ2� �LKK'	bV#�����)�~�/d2��a�0��_w�Y,YYY�$�cx�'��޸q�S����\�p��+����	�����!��p81�>    �����?������JEjg]ZZ�p����r��Q�B�V�B#�$I�<.� � ��x<�t�ZN��Ł@��ĩ��� �/��`p��#UUU:�6��(V8N��Dy|~�u(nh�"�HԽ�~Gg���M$%%�	����Ym�wt��|�h}��������[���ݺֶ�T�ۚ7o�F���la
#���m6��,�F��d�����I�L*�/_��n�[�/_�"�JE"�]��5�
>ER˫�W��NL�����$qVVoo_Eyy�����uZ-I����9:]$�|TR�6����[�l�t����@����x�'��l�#Cq��;n��0L$iko_�vmAA��ۜzc�c�h5���i��{oՊ���l�BQQQ����t�&;�   �='��D��.]�3!�	��9��2.���&v�S!cb��'v����[][�JQ���Ss�����b�~��(3syUf0�����utv��].�V��نپ���O��q�P`,PZZ���cwuw��:�c�#b�cL�98����7���C�g����{n����^y��ի�p���������3���hط�u�����-�8�L�U�������"�h�T8�������#Y"��P��i����lhh�(/�i�w�O�飋FB�z+uN0U^VVz����D���w�V��]]{��Q�N��e�Y^�:2HU�ɤv�������dI��h91�svoz�D��@0`6����O��h4N�3��F�>���D���6�p8��4|o�-G������o"dL   �������VS���j���r���,�
�
�)���D9q3��������~�_�ǎ9�N;�߿�޿�����e���|���kj����:|��B�Puu�R��-��y��[����d2izF�cdd�;�(��������J7��4����G��7<^o����@!���5���P%��d2�@ x��WB����9�L���d�D���3� ���䓻^}�_^�Ş�e�t��t�raaюG�syܻ�'b�㺭��vs9��̌���G�d��N!��hj�F�b����𰝦�3�����-�oi0�gg�L&�vG8<O&���n�����i�ϧT(ɤ�n������ⱸL&�*I$##N6���&�;$Ir�\�X,B��nO�q8l�׋�gg��[w����8\�R� I���d˳Y3L�    ������`p|*�i��P8��xh����*�rj�$M�>�/;;�����!�J�b��^/�b�	�v�#���L?��)
��Ҧ�8<<����^��T�\N'���j�w���t:���A$H�p%HB��dd��#�w?��!� ~����U���ޞ��$�_���B��.��jii��Ȭ�\�&oH")�;9�3���m�_���7�gg�\�bEMM�Lv�Z�oZ��c���&�0��C�׮YSTT     s����ozB�`��h4�#G�Z��T�~h�ٷž��s;��G\3]ohh`��%%�W׮���{     ��
���     �[�<�     �mĄ�A    ����     ̱��{�,���    IEND�B`�