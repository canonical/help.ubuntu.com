<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Aviseringar och aviseringslistan</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html.sv" title="Ditt skrivbord">Skrivbord</a> › <a class="trail" href="shell-overview.html.sv#desktop" title="Anpassa ditt skrivbord">Anpassa ditt skrivbord</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Aviseringar och aviseringslistan</span></h1></div>
<div class="region">
<div class="contents pagewide"></div>
<section id="what"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Vad är en avisering?</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Om ett program eller en systemkomponent vill få tag i din uppmärksamhet, kommer en avisering att visas längst upp på skärmen, eller på din låsskärm.</p>
<p class="p">Om du exempelvis får ett nytt chattmeddelande eller ett nytt e-postmeddelande så kommer du att få en avisering som informerar dig om detta. Chattaviseringar ges specialbehandling och representeras av de individuella kontakterna som skickade chattmeddelandena till dig.</p>
<p class="p">Andra aviseringar har valbara knappar. För att stänga en avisering av denna typ utan att välja en av dess alternativ, klicka på stängknappen.</p>
<p class="p">Att klicka på stängknappen på vissa aviseringar förkastar dem. Andra, som Rhythmbox eller ditt chattprogram kommer att förbli gömda i aviseringslistan.</p>
</div></div>
</div></section><section id="notificationlist"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Aviseringslistan</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Aviseringslistan ger dig ett sätt att få tillbaka dina aviseringar när det är bekvämt för dig. Den visas när du klickar på klockan eller trycker <span class="keyseq"><span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span>+<span class="key"><kbd>V</kbd></span></span>. Aviseringslistan innehåller alla aviseringar som du inte har agerat på eller som finns där permanent.</p>
<p class="p">Du kan visa en avisering genom att klicka på den i listan. Du kan stänga aviseringslistan genom att trycka <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>V</kbd></span></span> igen eller <span class="key"><kbd>Esc</kbd></span>.</p>
<p class="p">Klicka på knappen <span class="gui">Töm lista</span> för att tömma aviseringslistan.</p>
</div></div>
</div></section><section id="hidenotifications"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Dölja aviseringar</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Om du arbetar med något och inte vill bli störd kan du stänga av aviseringar.</p>
<p class="p">Du kan dölja alla aviseringar genom att öppna aviseringslistan och slå på <span class="gui">Stör ej</span> längst ner. Alternativt kan du:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Inställningar</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Inställningar</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Aviseringar</span> i sidopanelen för att öppna panelen.</p></li>
<li class="steps"><p class="p">Slå av <span class="gui">Stör ej</span>.</p></li>
</ol></div></div></div>
<p class="p">När de är avstängda kommer de flesta aviseringar inte att poppa upp längst upp på skärmen. Aviseringar kommer fortfarande att finnas tillgängliga i aviseringslistan när du visar den (genom att klicka på klockan, eller trycka på <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>V</kbd></span></span>) och de kommer att börja poppa upp igen när du slår på inställningen igen.</p>
<p class="p">Du kan också inaktivera eller återaktivera aviseringar för individuella program från panelen <span class="gui">Aviseringar</span>.</p>
</div></div>
</div></section><section id="lock-screen-notifications"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Dölja aviseringar på låsskärmen</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">När din skärm är låst, kommer aviseringar att visas på låsskärmen. Du kan av säkerhetsskäl konfigurera så att låsskärmen gömmer dessa aviseringar.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">För att slå av aviseringar när din skärm är låst:</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Inställningar</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Inställningar</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Aviseringar</span> i sidopanelen för att öppna panelen.</p></li>
<li class="steps"><p class="p">Slå av <span class="gui">Aviseringar på låsskärm</span>.</p></li>
</ol></div>
</div></div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html.sv#desktop" title="Anpassa ditt skrivbord">Anpassa ditt skrivbord</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
