<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Hitta en borttappad fil</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Hitta en borttappad fil</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du skapat eller hämtat en fil men inte kan hitta den, följ dessa tips.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Om du inte kommer ihåg var du sparade filen, men har en idé om vad du kallade den kan du <span class="link"><a href="files-search.html.sv" title="Sök efter filer">söka efter filen efter namn</a></span>.</p></li>
<li class="list"><p class="p">Om du nyss hämtade filen kan din webbläsare automatiskt ha sparat den till en gemensam mapp. Kontrollera mapparna <span class="file">Skrivbord</span> och <span class="file">Hämtningar</span> i din hemmapp.</p></li>
<li class="list"><p class="p">Du kan av misstag ha tagit bort filen. När du tar bort en fil flyttas den till papperskorgen där den stannar kvar tills du manuellt tömmer papperskorgen. Se <span class="link"><a href="files-recover.html.sv" title="Återskapa en fil från Papperskorgen">Återskapa en fil från Papperskorgen</a></span> för att lära dig hur du återställer en borttagen fil.</p></li>
<li class="list"><p class="p">Du kan ha bytt namn på filen på ett sätt som gjort filen dold. Filer som börjar med en <span class="file">.</span> eller slutar med ett <span class="file">~</span> är gömda för filhanteraren. Klicka på knappen visningsalternativ i verktygsfältet i <span class="app">Filer</span> och aktivera <span class="gui">Visa dolda filer</span> för att visa dem. Se <span class="link"><a href="files-hidden.html.sv" title="Dölj en fil">Dölj en fil</a></span> för att lära dig mer.</p></li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html.sv#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-recover.html.sv" title="Återskapa en fil från Papperskorgen">Återskapa en fil från Papperskorgen</a><span class="desc"> — Borttagna filer skickas normalt till Papperskorgen, men kan återställas.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
