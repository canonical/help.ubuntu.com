<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Låtar visas inte på min iPod när jag kopierar över dem</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Låtar visas inte på min iPod när jag kopierar över dem</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">När du kopplar en iPod till din dator kommer den att visas i ditt musikspelarprogram och också i filhanteraren (programmet <span class="app">Filer</span> i översiktsvyn <span class="gui">Aktiviteter</span>). Du måste kopiera låtar till din iPod via musikspelaren — om du kopierar dem via filhanteraren så kommer det inte att fungera eftersom låtarna inte kommer att hamna på rätt ställe. IPod:ar har en speciell plats för att spara låtar som musikspelarprogrammet känner till hur man når, men som filhanteraren inte känner till.</p>
<p class="p">Du måste också vänta på att låtarna ska sluta kopieras till iPod:en innan du kopplar från den. Innan du kopplar från iPod:en, försäkra dig om att du valt att göra en <span class="link"><a href="files-removedrive.html" title="Säker borttagning av extern enhet">säker borttagning av den</a></span>. Detta kommer att säkerställa att alla låtarna har kopierats korrekt.</p>
<p class="p">Ytterligare ett skäl till varför låtar kanske inte syns på din iPod kan vara att musikspelarprogrammet du använder inte har stöd för att konvertera låtarna från ett ljudformat till ett annat. Om du kopierar en låt som är sparade i ett ljudformat som inte har stöd för din iPod (till exempel en Ogg Vorbis-fil (.oga)) kommer musikspelaren att försöka konvertera den till ett format som iPod:en förstår, exempelvis MP3. Om det lämpliga konverteringsprogrammet (också känt som kodek eller kodare) inte är installerat kommer musikspelaren inte att kunna konvertera och kommer därför inte att kopiera låten. Leta i programinstalleraren efter en lämplig kodek.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
