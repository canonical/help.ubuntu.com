<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Jag kan inte höra några ljud alls från datorn</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="media.html#sound" title="Grundinställningar ljud">Ljud</a> » <a class="trail" href="sound-broken.html" title="Ljudproblem">Ljudproblem</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="sound-broken.html" title="Ljudproblem">Ljudproblem</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Jag kan inte höra några ljud alls från datorn</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Om du inte kan höra några ljud alls från din dator, till exempel när du försöker spela musik, prova dessa felsökningssteg för att se om du kan fixa problemet.</p></div>
<div id="mute" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Säkerställ att ljudvolymen inte är tyst</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Klicka på <span class="gui">ljudmenyn</span> i menyraden (den ser ut som en högtalare) och se till att ljudet inte är tystat eller satt till en låg volym.</p>
<p class="p">Vissa bärbara datorer har tangenter för att tysta ljudet på tangentbordet — tryck på den knappen för att se om det ljudet fungerar.</p>
<p class="p">Du bör också kontrollera att du inte har tystat programmet du använder för att spela upp ljud (t.ex. din musikspelare eller filmspelare). Programmet kan ha en tyst- eller volymknapp i dess huvudfönster, så kontrollera det också. Klicka också på ljudmenyn på menyraden och välj <span class="gui">Ljudinställningar</span>. När fönstret <span class="gui">Ljud</span> visas, gå till fliken <span class="gui">Program</span> och kontrollera att ditt program inte är tystat.</p>
</div></div>
</div></div>
<div id="speakers" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kontrollera att högtalarna är igång och korrekt anslutna</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Om din dator har externa högtalare, försäkra dig om att de är påslagna och att volymen är uppskruvad. Säkerställ att högtalarkabeln är ordentligt inkopplad i kontakten “ljudutgång“ på din dator. Denna kontakt är vanligtvis ljusgrön till färgen.</p>
<p class="p">Vissa ljudkort kan växla vilken kontakt som de använder som utgång (till högtalarna) och ingång (från till exempel en mikrofon). Utgångskontakten kan vara olika när du kör Linux än i Windows eller Mac OS. Prova att koppla in högtalarkabeln i olika ljudkontakter på datorn för att se om det fungerar.</p>
<p class="p">En sista sak att kontrollera är att se om ljudkabeln är ordentligt inkopplad på baksidan av högtalarna. Vissa högtalare har dessutom mer än en ingång.</p>
</div></div>
</div></div>
<div id="device" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kontrollera att rätt ljudenhet är vald</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Vissa datorer har flera “ljudenheter“ installerade. Vissa av dessa är kapabla att sända ut ljud medan andra inte är det, så du bör kontrollera att du har valt den rätta enheten. Det kan behövas ett antal försök för att hitta den rätta.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="gui">ljudmenyn</span> i <span class="gui">menyraden</span> och klicka på <span class="gui">Ljudinställningar</span>.</p></li>
<li class="steps"><p class="p">I fönstret <span class="gui">Ljud</span> som visas, testa en annan utmatning från listan <span class="gui">Spela ljud genom</span>.</p></li>
<li class="steps"><p class="p">För den valda enheten, klicka på <span class="gui">Testa ljud</span>. I fönstret som dyker upp, klicka på knappen för varje högtalare. Varje knapp kommer läsa upp sin position, bara i den kanal som motsvaras av den högtalaren.</p></li>
<li class="steps"><p class="p">Om det inte fungerar kan du behöva göra detsamma för de andra enheterna som är listade.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="hardware-detected" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kontrollera att ljudkortet detekterades ordentligt</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Ditt ljudkort kanske inte upptäcktes korrekt. I så fall kommer din dator tro att den inte kan spela upp ljud. En möjlig anledning till att kortet inte upptäcks korrekt är att drivrutinerna för kortet inte är installerade.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Gå till <span class="link"><a href="unity-dash-intro.html" title="Hitta program, filer, musik med mera med Snabbstartspanelen">Snabbstartspanelen</a></span> och öppna Terminalen.</p></li>
<li class="steps"><p class="p">Skriv <span class="cmd">aplay -l</span> och tryck <span class="key"><kbd>Retur</kbd></span>.</p></li>
<li class="steps"><p class="p">En lista över enheter kommer visas. Om det inte finns några <span class="gui">hårdvaruenheter för uppspelning</span> har ditt ljudkort inte upptäckts.</p></li>
</ol></div></div></div>
<p class="p">Om ditt ljudkort inte upptäckts kan du behöva installera drivrutinerna manuellt. Hur det går till beror på vilket kort du har.</p>
<p class="p">Du kan se vilket ljudkort du har genom att använda kommandot <span class="cmd">lspci</span> i <span class="app">Terminalen</span>. Du får ett mer fullständigt resultat om du kör <span class="cmd">lspci</span> som <span class="link"><a href="user-admin-explain.html" title="Hur fungerar administratörsbehörighet?">superanvändare</a></span>; skriv <span class="cmd">sudo lspci</span> och skriv ditt lösenord. Se om en <span class="em">ljudkontroll</span> eller <span class="em">ljudenhet</span> visas i listan—den bör visa ljudkortets tillverkare och modellnummer. <span class="cmd">sudo lspci -v</span> visar en lista med mer detaljerad information.</p>
<p class="p">Du kan hitta och installera drivrutiner för ditt kort genom att söka på internet. Annars kan du <span class="link"><a href="report-ubuntu-bug.html" title="Rapportera ett problem i Ubuntu">göra en felanmälan</a></span>.</p>
<p class="p">Om du inte kan få tag i drivrutiner för ditt ljudkort kanske du föredrar att köpa ett nytt ljudkort. Du kan köpa ljudkort som kan installeras inuti dator eller externa USB-ljudkort.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="sound-broken.html" title="Ljudproblem">Ljudproblem</a><span class="desc"> — Felsök problem som att inte få ljud eller få dåligt ljudkvalitet.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
