<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>pam_motd</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="other-useful-applications.html" title="Ytterligare användbara program">Ytterligare användbara program</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="other-useful-applications.html" title="Ytterligare användbara program">Föregående</a><a class="nextlinks-next" href="etckeeper.html" title="etckeeper">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">pam_motd</h1></div>
<div class="region">
<div class="contents">
<p class="para">När du loggat in till en Ubuntu server så har du kanske sätt det informativa Message Of The Day (MOTD). Denna information inhämtas och visas genom att använda några paket:</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
        <p class="para">
        <span class="em emphasis">landscape-common:</span> provides the core libraries of <span class="app application">landscape-client</span>,
	which is needed to manage systems with <a href="http://landscape.canonical.com/" class="ulink" title="http://landscape.canonical.com/">Landscape</a> (proprietary).  Yet the package also includes
        the <span class="app application">landscape-sysinfo</span> utility which is responsible for displaying core system data involving cpu, memory, disk space, etc.  For instance:
        </p>

<div class="screen"><pre class="contents "><span class="output computeroutput">
	  System load:  0.0               Processes:           76
	  Usage of /:   30.2% of 3.11GB   Users logged in:     1
	  Memory usage: 20%               IP address for eth0: 10.153.107.115
	  Swap usage:   0%

	  Graph this data and manage this system at https://landscape.canonical.com/
</span>
</pre></div>

        <div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
                <p class="para">
                You can run landscape-sysinfo manually at any time.
                </p>
        </div></div></div></div>

      </li>
<li class="list itemizedlist">
        <p class="para">
        <span class="em emphasis">update-notifier-common:</span> provides information on available package updates, impending filesystem checks (fsck), and required reboots (e.g.: after a kernel upgrade).
        </p>
      </li>
</ul></div>
<p class="para">    
    <span class="app application">pam_motd</span> executes the scripts in <span class="file filename">/etc/update-motd.d</span> in order based on the number 
    prepended to the script.  The output of the scripts is written to <span class="file filename">/var/run/motd</span>, keeping the numerical order, 
    then concatenated with <span class="file filename">/etc/motd.tail</span>.
    </p>
<p class="para">Du kan lägga till din egna dynamiska information till MOTD. Till exempel, för att lägga till lokal väderinformation:</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
        <p class="para">Installera först paketet <span class="app application">weather-util</span>:</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo apt-get install weather-util</span>
</pre></div>

      </li>
<li class="list itemizedlist">
        <p class="para">Verktyget <span class="app application">weather</span> använder METAR-data från National Oceanic and Atmospheric Administration och prognoser från National Weather Service. För att hitta lokal information behöver du ICAO platsindikator på 4 tecken. Den kan du ta reda på genom att bläddra i webbplatsen <a href="http://www.weather.gov/tg/siteloc.shtml" class="ulink" title="http://www.weather.gov/tg/siteloc.shtml">National Weather Service</a>.</p>

        <p class="para">Även om National Weather Service är en amerikansk myndighet finns det väderstationer över hela världen. Men det lokala vädret för alla platser utanför USA kanske inte är tillgängliga.</p>
      </li>
<li class="list itemizedlist">
        <p class="para">Skapa <span class="file filename">/usr/local/bin/local-weather</span>, ett enkelt skal-skript till att använda <span class="app application">weather</span> med din lokala ICAO-indikator:</p>

<div class="code"><pre class="contents ">#!/bin/sh
#
#
# Prints the local weather information for the MOTD.
#
#

# Replace KINT with your local weather station.
# Local stations can be found here: http://www.weather.gov/tg/siteloc.shtml

echo
weather -i KINT
echo

</pre></div>
      </li>
<li class="list itemizedlist">
        <p class="para">Gör skriptet exekverbart:</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo chmod 755 /usr/local/bin/local-weather</span>
</pre></div>
      </li>
<li class="list itemizedlist">
        <p class="para">
        Next, create a symlink to <span class="file filename">/etc/update-motd.d/98-local-weather</span>:
        </p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo ln -s /usr/local/bin/local-weather /etc/update-motd.d/98-local-weather</span>
</pre></div>
      </li>
<li class="list itemizedlist">
        <p class="para">
        Finally, exit the server and re-login to view the new MOTD.
        </p>
      </li>
</ul></div>
<p class="para">
    You should now be greeted with some useful information, and some information about the local weather that may not be
    quite so useful. Hopefully the <span class="app application">local-weather</span> example demonstrates the flexibility of
    <span class="app application">pam_motd</span>.
    </p>
</div>
<div class="links sectionlinks" role="navigation"><ul><li class="links"><a class="xref" href="pam_motd.html#pam_motd-resources" title="Resurser">Resurser</a></li></ul></div>
<div class="sect2 sect" id="pam_motd-resources"><div class="inner">
<div class="hgroup"><h2 class="title">Resurser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
	<p class="para">
        See the <a href="http://manpages.ubuntu.com/manpages/trusty/en/man5/update-motd.5.html" class="ulink" title="http://manpages.ubuntu.com/manpages/trusty/en/man5/update-motd.5.html">update-motd man page</a> for
        more options available to <span class="app application">update-motd</span>.
	</p>
	</li>
<li class="list itemizedlist">
        <p class="para">Debian Package of the Day har en <a href="http://debaday.debian.net/2007/10/04/weather-check-weather-conditions-and-forecasts-on-the-command-line/" class="ulink" title="http://debaday.debian.net/2007/10/04/weather-check-weather-conditions-and-forecasts-on-the-command-line/">väder</a>-artikel som har mer detaljer om att använda verktyget <span class="app application">weather</span>.</p>
        </li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="other-useful-applications.html" title="Ytterligare användbara program">Föregående</a><a class="nextlinks-next" href="etckeeper.html" title="etckeeper">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
