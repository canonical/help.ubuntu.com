<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Säkerhet &amp; sekretess</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Säkerhet &amp; sekretess</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Den här sidan beskriver inställningarna i modulen <span class="app">Säkerhet &amp; sekretess</span>. Fönstret har fyra flikar:</p></div>
<div id="tab1" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Säkerhet</span></h2></div>
<div class="region"><div class="contents"><p class="p">Dessa inställningar anger huruvida ett lösenord behöver anges när Ubuntu vaknar upp från <span class="link"><a href="power-suspend.html" title="Vad händer när jag försätter min dator i vänteläge?">vänteläge</a></span> eller för att återvända från en blank skärm. Din dator blir säkrare om lösenord krävs i de fallen.</p></div></div>
</div></div>
<div id="tab2" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Filer &amp; Program</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Dessa inställningar låter dig ange vilka av senast använda filer, mappar och program som listas i t ex <span class="gui">Dash</span>.</p>
<p class="p">För att bestämma senast använda filer, mappar och program, samlar Ubuntu in användningsdata. Om du önskar, kan du stänga <span class="gui">AV</span> insamling av användningsdata och rensa bort en del eller all insamlad användningsdata.</p>
<p class="p"><span class="gui">Inkludera:</span>-listan tar upp några vanliga filtyper. För att inkludera en filtyp i användningsdatan, markera boxen näst intill. För att exkludera en filtyp från användningsdatan, avmarkera motsvarande box.</p>
<p class="p"><span class="gui">Uteslut:</span>-listan anger mappar och program som exkluderas från användningsdatan. För att lägga till en mapp eller program till listan, klicka på "+"-knappen och välj en mapp eller ett program. För att ta bort en mapp eller program från listan, markera mappen eller programmet och klicka på "-"-knappen.</p>
</div></div>
</div></div>
<div id="tab3" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Sök</span></h2></div>
<div class="region"><div class="contents"><p class="p">Den här inställningen anger huruvida sökresultat från internet skall inkluderas vid sökning i <span class="gui">Dash</span>. För mer information om sökresultat från internet, och företagen som tillhandahåller dem, se Canonicals sekretesspolicy som du kan nå från <span class="gui">Diagnostik</span>-fliken.</p></div></div>
</div></div>
<div id="tab4" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Diagnostik</span></h2></div>
<div class="region"><div class="contents"><p class="p">Dessa inställningar anger vilken typ av systeminformation som Ubuntu kan skicka till Canonical. Informationen (om du tillåter att den skickas) hjälper Canonical att förbättra Ubuntu. Om du vill veta mer om hur Canonical använder systeminformationen, klicka på <span class="gui">Sekretesspolicy</span> för att läsa Canonicals sekretesspolicy.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html" title="Användarkonton">användarkonton</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="display-lock.html" title="Lås automatiskt din skärm">Lås automatiskt din skärm</a><span class="desc"> — Hindra andra från att använda ditt skrivbord när du lämnar datorn.</span>
</li>
<li class="links ">
<a href="net-security-tips.html" title="Trygghet på internet">Trygghet på internet</a><span class="desc"> — Allmänna tips när du använder internet</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
