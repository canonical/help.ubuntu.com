<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ta bort filer och mappar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Ta bort filer och mappar</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du inte längre vill ha en fil eller mapp kan du ta bort den. När du tar bort något flyttas det till <span class="gui">Papperskorgen</span>, där det förvaras tills du tömmer papperskorgen. Du kan <span class="link"><a href="files-recover.html" title="Återställ en fil från Papperskorgen">återställa objekten</a></span> i <span class="gui">Papperskorgen</span> till deras ursprungliga plats om du vill ha tillbaka dem, eller om de togs bort av misstag.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">För att skicka en fil till papperskorgen:</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Välj objektet du vill placera i papperskorgen genom att klicka på det en enda gång.</p></li>
<li class="steps"><p class="p">Tryck <span class="key"><kbd>Delete</kbd></span> på ditt tangentbord. Du kan också dra objektet till <span class="gui">Papperskorgen</span> i sidoraden.</p></li>
</ol></div>
</div></div>
<p class="p">För att ta bort filer permanent, och frigöra diskutrymme på din dator, måste du tömma papperskorgen. För att tömma papperskorgen, högerklicka på <span class="gui">Papperskorgen</span> i sidoraden och välj <span class="gui">Töm papperskorgen</span>.</p>
</div>
<div id="permanent" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ta bort en fil permanent</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan ta bort en fil permanent direkt, utan att först behöva skicka den till papperskorgen.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">För att ta bort en fil permanent:</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Markera objektet som du vill ta bort.</p></li>
<li class="steps"><p class="p">Håll ner <span class="key"><kbd>Shift</kbd></span>-tangenten, och tryck sedan på <span class="key"><kbd>Delete</kbd></span>-tangenten på ditt tangentbord.</p></li>
<li class="steps"><p class="p">Eftersom du inte kan ångra det här kommer du få bekräfta att du verkligen vill ta bort filen eller mappen.</p></li>
</ol></div>
</div></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du ofta behöver ta bort filer utan att använda papperskorgen (om du till exempel ofta arbetar med känslig information) kan du lägga till en <span class="gui">Ta bort</span>-post i högerklickmenyn för filer och mappar. Klicka på <span class="gui">Filer</span> i menyraden, välj <span class="gui">Inställningar</span> och välj fliken <span class="gui">Beteende</span>. Välj <span class="gui">Inkludera ett Ta bort-kommando som förbigår Papperskorgen</span>.</p></div></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Raderade filer på en <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">flyttbar enhet</a></span> kanske inte syns i andra operativsystem, som Windows eller Mac OS. Filerna finns kvar, och kommer bli tillgängliga när du ansluter enheten igen.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="nautilus-behavior.html#trash" title="Papperskorg">Filhanterarens papperskorginställningar</a></li>
<li class="links ">
<a href="files-recover.html" title="Återställ en fil från Papperskorgen">Återställ en fil från Papperskorgen</a><span class="desc"> — Borttagna filer skickas normalt till Papperskorgen, men kan återställas.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
