<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Välj ditt lösenord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="user-accounts.html" title="Användarkonton">Användare</a> › <a class="trail" href="user-accounts.html#passwords" title="Lösenord">Lösenord</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Välj ditt lösenord</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Det är en bra idé att byta lösenord med jämna mellanrum, särskilt om du tror att någon annan känner till ditt lösenord.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ikonen längst till höger i <span class="gui">menylisten</span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Öppna <span class="gui">Användarkonton</span>.</p></li>
<li class="steps">
<p class="p">Klicka på etiketten bredvid <span class="gui">Lösenord</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Etiketten bör se ut som en serie prickar eller rutor om du redan har ett lösenord.</p></div></div></div></div>
</li>
<li class="steps">
<p class="p">Skriv in ditt nuvarande lösenord, och skriv sedan in det nya lösenordet. Skriv ditt nya lösenord igen i fältet <span class="gui">Bekräfta lösenord</span>.</p>
<p class="p">Du kan också klicka på knappen bredvid fältet <span class="gui">Nytt lösenord</span> för att välja ett slumpgenererat säkert lösenord. Dessa lösenord är svåra för andra att gissa sig fram till, men de kan vara svåra att lägga på minnet, så var försiktig.</p>
</li>
<li class="steps"><p class="p">Klicka på <span class="gui">Ändra</span>.</p></li>
</ol></div></div></div>
<p class="p">Var noga med att <span class="link"><a href="user-goodpassword.html" title="Välj ett säkert lösenord">välja ett bra lösenord</a></span>. Detta hjälper dig skydda ditt användarkonto.</p>
</div>
<div id="changepass" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ändra nyckelknippans lösenord</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Om du ändrar inloggningslösenord kan det tappa synkronisering med <span class="em">nyckelknippans lösenord</span>. Nyckelknippan gör att du inte behöver komma ihåg många olika lösenord genom att bara kräva ett <span class="em">master-lösenord</span> för att komma åt allihop. Om du ändrar ditt användarlösenord (se ovan) kommer ditt lösenord till nyckelknippan vara samma som ditt gamla lösenord. För att ändra nyckelknippans lösenord (för att stämma överens med ditt inloggningslösenord):</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna programmet <span class="app">Lösenord och nycklar</span> från <span class="gui">Snabbstartspanelen</span>.</p></li>
<li class="steps"><p class="p">I menyn <span class="gui">Visa</span>, kontrollera att <span class="gui">Enligt nyckelknippa</span> är markerad.</p></li>
<li class="steps"><p class="p">I sidpanelen under <span class="gui">Lösenord</span>, högerklicka på <span class="gui">Inloggningsnyckelknippa</span> och välj <span class="gui">Byt lösenord</span>.</p></li>
<li class="steps"><p class="p">Skriv in <span class="gui">Gammalt lösenord</span>, följt av ditt nya <span class="gui">Lösenord</span>, och <span class="gui">Bekräfta</span> ditt nya lösenord genom att skriva in det igen.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">OK</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="user-accounts.html#passwords" title="Lösenord">Lösenord</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="user-goodpassword.html" title="Välj ett säkert lösenord">Välj ett säkert lösenord</a><span class="desc"> — Använd längre och mer komplicerade lösenord.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
