<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Virtualisering</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = "index.html.en";
        } else {
                window.location = href.replace(/\.html.*/, ".html.en");
        }
         return false;
      }
      function browserPreferredLanguage() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = href;
        } else {
                window.location = href.replace(/\.html.*/, ".html");
        }
        return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../18.04" class="trail">Ubuntu 18.04</a> » <a class="trail" href="index.html.sv" title="Ubuntu serverguide">Ubuntu serverguide</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="bacula.html.sv" title="Bacula">Föregående</a><a class="nextlinks-next" href="libvirt.html.sv" title="libvirt">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Virtualisering</h1></div>
<div class="region">
<div class="contents">
<p class="para">Virtualisering används i många olika miljöer och situationer. Om du är en utvecklare så kan virtualisering tillhandahålla en begränsad miljö där du på ett säkert sätt utföra nästan alla typer av utveckling utan risk att förstöra din huvudsakliga arbetsmiljö. Om du är en systemadministratör så kan du använda virtualisering för att enklare separera dina tjänster och på förfrågan flytta dem.</p>
<p class="para">The default virtualization technology supported in Ubuntu is
  <span class="app application">KVM</span>. For Intel and AMD hardware KVM requires
  virtualization extensions. But KVM is also available for IBM Z and LinuxONE,
  IBM POWER as well as for ARM64.
  <span class="app application">Xen</span> is also supported on Ubuntu, but not for all architecture, 
  for example not for IBM Z and LinuxONE.
  Xen can take advantage of virtualization extensions,
  when available, but can also be used on hardware without virtualization
  extensions. <span class="app application">Qemu</span> is another popular solution for
  hardware without virtualization extensions.</p>
</div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="libvirt.html.sv" title="libvirt">libvirt</a></li>
<li class="links"><a class="xref" href="qemu.html.sv" title="Qemu">Qemu</a></li>
<li class="links"><a class="xref" href="cloud-images-and-uvtool.html.sv" title="Cloud images and uvtool">Cloud images and uvtool</a></li>
<li class="links"><a class="xref" href="ubuntucloud.html.sv" title="Ubuntu Cloud">Ubuntu Cloud</a></li>
<li class="links"><a class="xref" href="lxd.html.sv" title="LXD">LXD</a></li>
<li class="links"><a class="xref" href="lxc.html.sv" title="LXC">LXC</a></li>
</ul></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="bacula.html.sv" title="Bacula">Föregående</a><a class="nextlinks-next" href="libvirt.html.sv" title="libvirt">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address
          so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>
          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p>
</div>
</div>
</body>
</html>
