<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Maskinvara och drivrutiner</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Maskinvara och drivrutiner</span></h1></div>
<div class="region">
<div class="contents">
<div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-grid ">
<div class="links-grid-link"><a href="bluetooth.html" title="Bluetooth">Bluetooth</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="bluetooth-connect-device.html" title="Anslut din dator till en Bluetooth-enhet">Anslut</a></span>, <span class="link"><a href="bluetooth-send-file.html" title="Skicka filer till en Bluetooth-enhet">skicka filer</a></span>, <span class="link"><a href="bluetooth-turn-on-off.html" title="Aktivera eller inaktivera Bluetooth">aktivera och inaktivera</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="disk.html" title="Diskar och lagring">Diskar och lagring</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="disk-capacity.html" title="Kontrollera hur mycket diskutrymme som finns kvar">Diskutrymme</a></span>, <span class="link"><a href="disk-benchmark.html" title="Testa din hårddisks prestanda">prestanda</a></span>, <span class="link"><a href="disk-check.html" title="Kontrollera din hårddisk efter problem">problem</a></span>, <span class="link"><a href="disk-partitions.html" title="Hantera volymer och partitioner">volymer och partitioner</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="hardware-auth.html" title="Fingeravtryck &amp; smartkort">Fingeravtryck &amp; smartkort</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="session-fingerprint.html" title="Logga in med ett fingeravtryck">Fingeravtrycksläsare</a></span>, smartkort…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="color.html" title="Färghantering">Färghantering</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="color-whyimportant.html" title="Varför är färghantering viktigt?">Varför är detta viktigt</a></span>, <span class="link"><a href="color.html#profiles" title="Färgprofiler">Färgprofiler</a></span>, <span class="link"><a href="color.html#calibration" title="Kalibrering">Hur du kalibrerar en enhet</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="mouse.html" title="Mus">Mus</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="mouse-lefthanded.html" title="Använd din mus med vänster hand">Vänsterhänt</a></span>, <span class="link"><a href="mouse-sensitivity.html" title="Justera hastigheten för musen och styrplattan">hastighet och känslighet</a></span>, <span class="link"><a href="mouse-touchpad-click.html" title="Klicka, dra eller rulla med styrplattan">klickning och rullning med styrplatta</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="power.html" title="Ström och batteri">Ström och batteri</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="power-status.html" title="Kontrollera batteristatus">Batteristatus</a></span>, <span class="link"><a href="power-suspend.html" title="Vad händer när jag försätter min dator i vänteläge?">försätta i vänteläge</a></span>, <span class="link"><a href="power-whydim.html" title="Varför tonas min skärm ner efter ett tag?">skärmtoning</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="keyboard-layouts.html" title="Använd alternativa tangentbordslayouter">Tangentbordslayouter</a></span>, <span class="link"><a href="keyboard-cursor-blink.html" title="Få tangentbordsmarkören att blinka">markörblinkning</a></span>, <span class="link"><a href="a11y.html#mobility" title="Rörelsehinder">tangentbordshjälpmedel</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="printing.html" title="Utskrifter">Utskrifter</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="printing-setup.html" title="Ställ in en lokal skrivare">Lokal inställning</a></span>, <span class="link"><a href="printing-order.html" title="Skriv ut sidor i en annan ordning">ordna och sortera</a></span>, <span class="link"><a href="printing-2sided.html" title="Skriv ut dubbelsidigt och flersidslayouter">dubbelsidig och flersidig utskrift</a></span>…</span></div>
</div>
</div></div></div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Fler ämnen</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="hardware-driver.html" title="Vad är en drivrutin?">Vad är en drivrutin?</a><span class="desc"> — En hårdvaru-/enhetsdrivrutin låter din dator använda enheter som ansluts till den.</span>
</li></ul></div>
</div></div>
</div>
<div id="problems" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Vanliga problem</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region"><ul>
<li class="links "><a href="bluetooth.html#problems" title="Problem">Bluetooth-problem</a></li>
<li class="links ">
<a href="net-wireless-troubleshooting.html" title="Felsökning av trådlösa nätverk">Felsökning av trådlösa nätverk</a><span class="desc"> — Identifiera och fixa problem med trådlösa anslutningar.</span>
</li>
<li class="links ">
<a href="sound-broken.html" title="Ljudproblem">Ljudproblem</a><span class="desc"> — Felsök problem som att inte få ljud eller få dåligt ljudkvalitet.</span>
</li>
<li class="links ">
<a href="hardware-cardreader.html" title="Problem med mediakortsläsare">Problem med mediakortsläsare</a><span class="desc"> — Felsök mediakortsläsare</span>
</li>
<li class="links ">
<a href="printing.html#problems" title="Skrivarproblem">Skrivarproblem</a><span class="desc"> — Skrivare som inte detekterats, papper som fastnat, utskrifter som ser fel ut…</span>
</li>
<li class="links ">
<a href="hardware-problems-graphics.html" title="Skärmproblem">Skärmproblem</a><span class="desc"> — Felsök skärm- och grafikproblem.</span>
</li>
<li class="links ">
<a href="power.html#problems" title="Problem">Strömproblem</a><span class="desc"> — Felsök problem med ström och batterier.</span>
</li>
</ul></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
