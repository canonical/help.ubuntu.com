<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Visning och skärm</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Visning och skärm</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="display-dual-monitors.html" title="Anslut en extern skärm till din bärbara dator"><span class="title">Anslut en extern skärm till din bärbara dator</span><span class="linkdiv-dash"> — </span><span class="desc">Använd två skärmar för din bärbara dator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="display-dual-monitors-desktop.html" title="Anslut en extraskärm"><span class="title">Anslut en extraskärm</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in två skärmar för din skrivbordsdator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="look-background.html" title="Byt skrivbordsbakgrund"><span class="title">Byt skrivbordsbakgrund</span><span class="linkdiv-dash"> — </span><span class="desc">Ange en bild, färg, eller färgskala som skrivbordsbakgrund.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="display-lock.html" title="Lås automatiskt din skärm"><span class="title">Lås automatiskt din skärm</span><span class="linkdiv-dash"> — </span><span class="desc">Hindra andra från att använda ditt skrivbord när du lämnar datorn.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="session-screenlocks.html" title="Skärmen låser sig själv allt för snabbt"><span class="title">Skärmen låser sig själv allt för snabbt</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra hur lång tid det får gå innan skärmen låses i inställningarna för <span class="gui">Ljusstyrka &amp; Lås</span>.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="display-dimscreen.html" title="Ställ in skärmens ljusstyrka"><span class="title">Ställ in skärmens ljusstyrka</span><span class="linkdiv-dash"> — </span><span class="desc">Minska skärmens ljusstyrka för att spara energi, eller öka ljusstyrkan för att göra den mer lättläst i starkt ljus.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="look-resolution.html" title="Ändra storlek och rotation för skärmen"><span class="title">Ändra storlek och rotation för skärmen</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra skärmens upplösning och dess orientering (rotation).</span></a></div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html" title="Användarkonton">användarkonton</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
