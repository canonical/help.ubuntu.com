<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skärmbilder och skärminspelningar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 20.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="tips.html.sv" title="Tips och tricks">Tips och tricks</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Skärmbilder och skärminspelningar</span></h1></div>
<div class="region">
<div class="contents pagewide"><p class="p">Du kan ta en bild av din skärm (en <span class="em">skärmbild</span>) eller spela in en video av vad som händer på skärmen (en <span class="em">skärminspelning</span>). Detta är användbart om du vill visa någon hur något görs på datorn, till exempel. Skärmbilder och skärminspelningar är normala bild- och videofiler, så du kan e-posta dem och dela dem på nätet.</p></div>
<section id="screenshot"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Ta en skärmbild</span></h2></div>
<div class="region">
<div class="contents pagewide"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna <span class="app">Skärmbild</span> från översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span>.</p></li>
<li class="steps"><p class="p">I fönstret <span class="app">Skärmbild</span>, välj huruvida hela skärmen, det aktuella fönstret eller ett område på skärmen ska avbildas. Sätt en fördröjning om du behöver välja ett fönster eller på annat sätt arrangera skrivbordet för skärmbilden. Välj sedan effekterna du vill ha.</p></li>
<li class="steps">
<p class="p">Klicka på <span class="gui">Ta skärmbild</span>.</p>
<p class="p">Om du valde <span class="gui">Välj området att fånga</span> kommer markören att ändras till ett hårkors. Klicka och dra ett område som du önskar avbilda.</p>
</li>
<li class="steps">
<p class="p">I fönstret <span class="gui">Spara skärmbild</span>, mata in ett filnamn och välj en mapp, klicka sedan på <span class="gui">Spara</span>.</p>
<p class="p">Alternativt, importera skärmbilden direkt i ett bildredigeringsprogram utan att spara det först. Klicka på <span class="gui">Kopiera till urklipp</span> och klistra sedan in bilden i det andra programmet eller dra miniatyrskärmbilden till programmet.</p>
</li>
</ol></div></div></div></div>
<section id="keyboard-shortcuts"><div class="inner">
<div class="hgroup pagewide"><h3 class="title"><span class="title">Tangentbordsgenvägar</span></h3></div>
<div class="region"><div class="contents pagewide">
<p class="p">Ta snabbt en skärmbild av skrivbordet, ett fönster eller ett område när som helst via dessa globala tangentbordsgenvägar:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="key"><kbd>Prt Scrn</kbd></span> för att ta en skärmbild av skrivbordet.</p></li>
<li class="list"><p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>uppåtpil</kbd></span></span> för att ta en skärmbild av ett fönster.</p></li>
<li class="list"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Prt Scrn</kbd></span></span> för att ta en skärmbild av ett område som du väljer.</p></li>
</ul></div></div></div>
<p class="p">När du använder en tangentbordsgenväg kommer bilden automatiskt att sparas i din mapp <span class="file">Bilder</span> med ett filnamn som börjar med <span class="file">Skärmbild</span> och inkluderar datum och tid då den togs.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Om du inte har en mapp <span class="file">Bilder</span>, kommer bilderna att sparas i din hemmapp istället.</p></div></div></div>
</div>
<p class="p">Du kan också hålla ner <span class="key"><kbd>Ctrl</kbd></span> med någon av ovanstående genvägar för att kopiera skärmbilden till urklipp istället för att spara den.</p>
</div></div>
</div></section>
</div>
</div></section><section id="screencast"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Gör en skärminspelning</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Du kan göra en videoinspelning av vad som händer på din skärm:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps">
<p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>R</kbd></span></span> för att börja spela in det som finns på din skärm.</p>
<p class="p">En röd cirkel visas i övre högra hörnet av skärmen när inspelningen pågår.</p>
</li>
<li class="steps"><p class="p">När du är klar tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>R</kbd></span></span> igen för att avsluta inspelningen.</p></li>
<li class="steps"><p class="p">Videon sparas automatiskt i din mapp <span class="file">Videor</span> med ett filnamn som börjar med <span class="file">Skärminspelning</span> och inkluderar datum och tid när den spelades in.</p></li>
</ol></div></div></div>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Om du inte har en mapp <span class="file">Videor</span>, kommer videorna att sparas i din hemmapp istället.</p></div></div></div>
</div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="tips.html.sv" title="Tips och tricks">Tips och tricks</a><span class="desc"> — <span class="link"><a href="tips-specialchars.html.sv" title="Mata in speciella tecken">Specialtecken</a></span>, <span class="link"><a href="mouse-middleclick.html.sv" title="Mittenklick">genvägar för mittenklick</a></span>…</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
