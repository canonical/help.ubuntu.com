<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Muspekaren rör sig inte</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 22.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus</a> › <a class="trail" href="mouse.html.sv#problems" title="Vanliga problem">Vanliga problem</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 22.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus</a> › <a class="trail" href="mouse.html.sv#problems" title="Vanliga problem">Vanliga problem</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Muspekaren rör sig inte</span></h1></div>
<div class="region">
<div class="contents pagewide"><div role="navigation" class="links sectionlinks"><div class="inner"><div class="region"><ul>
<li class="links "><a href="mouse-problem-notmoving.html.sv#plugged-in" title="Kontrollera att musen är ansluten">Kontrollera att musen är ansluten</a></li>
<li class="links "><a href="mouse-problem-notmoving.html.sv#broken" title="Kontrollera att musen verkligen fungerar">Kontrollera att musen verkligen fungerar</a></li>
<li class="links "><a href="mouse-problem-notmoving.html.sv#wireless-mice" title="Kontrollera trådlösa möss">Kontrollera trådlösa möss</a></li>
</ul></div></div></div></div>
<section id="plugged-in"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Kontrollera att musen är ansluten</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Om du har en mus med en kabel, kontrollera att den är ordentligt ansluten till din dator.</p>
<p class="p">Om det är en USB-mus (med en fyrkantig kontakt), prova att ansluta den till en annan USB-kontakt. Om det är en PS/2-mus (med en liten rund kontakt med sex stift), säkerställ att den anslutits till den gröna muskontakten snarare än den lila tangentbordskontakten. Du kan bli tvungen att starta om datorn om den inte var ansluten.</p>
</div></div>
</div></section><section id="broken"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Kontrollera att musen verkligen fungerar</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Anslut musen till en annan dator och se om den fungerar.</p>
<p class="p">Om musen är en optisk- eller lasermus bör ljus skina ut från musens undersida om den är påslagen. Om det inte finns något ljus, kontrollera att den är påslagen. Om den är det och det fortfarande inte finns något ljus kan musen vara trasig.</p>
</div></div>
</div></section><section id="wireless-mice"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Kontrollera trådlösa möss</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Säkerställ att musen är påslagen. Det finns ofta en knapp på undersidan av musen som slår av musen helt så att du kan ta den med dig utan att den vaknar upp hela tiden.</p></li>
<li class="list"><p class="p">Om du använder en Bluetooth-mus, försäkra dig om att du verkligen har parat ihop musen med din dator. Se <span class="link"><a href="bluetooth-connect-device.html.sv" title="Anslut din dator till en Bluetooth-enhet">Anslut din dator till en Bluetooth-enhet</a></span>.</p></li>
<li class="list"><p class="p">Klicka med en knapp och se om muspekaren flyttar sig nu. Vissa trådlösa möss kan försättas i strömsparläge för att spara ström, så de kan sluta svara tills du klicka med en knapp. Se <span class="link"><a href="mouse-wakeup.html.sv" title="Musen reagerar med fördröjning innan den börjar fungera">Musen reagerar med fördröjning innan den börjar fungera</a></span>.</p></li>
<li class="list"><p class="p">Kontrollera att musens batteri är laddat.</p></li>
<li class="list"><p class="p">Säkerställ att mottagaren (adapter) är ordentligt ansluten till datorn.</p></li>
<li class="list"><p class="p">Om din mus och mottagare kan användas på olika radiokanaler, kontrollera att båda är inställda på samma kanal.</p></li>
<li class="list"><p class="p">Du kan vara tvungen att trycka på en knapp på musen, mottagaren eller båda för att etablera en anslutning. Instruktionshandboken för din mus bör ha fler detaljer om detta är fallet.</p></li>
</ul></div></div></div>
<p class="p">De flesta trådlösa möss (radio) bör fungera automatiskt när du ansluter dem till din dator. Om du har en Bluetooth- eller IR-mus (Infraröd) kan du behöva genomföra några extra steg för att få den att fungera. Stegen kan bero på tillverkare och modell av din mus.</p>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="mouse.html.sv#problems" title="Vanliga problem">Vanliga musproblem</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
