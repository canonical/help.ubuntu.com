<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Share your desktop</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="sharing.html" title="Sharing">Sharing</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Share your desktop</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">You can let other people view and control your desktop from another computer
 with a desktop viewing application. Configure <span class="app">Desktop Sharing</span> to
 allow others to access your desktop and set the security preferences.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">In the <span class="gui">Dash</span>, open <span class="app">Desktop Sharing</span>.</p></li>
<li class="steps"><p class="p">To let others view your desktop, select
 <span class="gui">Allow other users to view your desktop</span>. This means that other
 people will be able to attempt to connect to your computer and view what's
 on your screen.</p></li>
<li class="steps"><p class="p">To let others interact with your desktop, select
 <span class="gui">Allow other users to control your desktop</span>. This may allow the
 other person to move your mouse, run applications, and browse files
 on your computer, depending on the security settings which you are currently
 using.</p></li>
</ol></div></div></div>
</div>
<div id="security" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Security</span></h2></div>
<div class="region"><div class="contents">
<p class="p">It is important that you consider the full extent of what each security
 option means before changing it.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Confirm access to your machine</dt>
<dd class="terms">
<p class="p">If you want to be able to choose whether to allow someone to access
 your desktop, select <span class="gui">You must confirm each access to this machine</span>.
 If you disable this option, you will not be asked whether you want to allow
 someone to connect to your computer.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">This option is enabled by default.</p></div></div></div></div>
</dd>
<dt class="terms">Enable password</dt>
<dd class="terms">
<p class="p">To require other people to use a password when connecting to your
 desktop, select <span class="gui">Require the user to enter this password</span>. If you do
 not use this option, anyone can attempt to view your desktop.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">This option is disabled by default, but you should enable it and set
 a secure password.</p></div></div></div></div>
</dd>
<dt class="terms">Allow access to your desktop over the Internet</dt>
<dd class="terms">
<p class="p">If your router supports UPnP Internet Gateway Device Protocol and it is
 enabled, you can allow other people who are not on your local network to view
 your desktop. To allow this, select <span class="gui">Automatically configure UPnP router to
 open and forward ports</span>. Alternatively, you can configure your router
 manually.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">This option is disabled by default.</p></div></div></div></div>
</dd>
</dl></div></div></div>
</div></div>
</div></div>
<div id="notification-icon" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Show notification area icon</span></h2></div>
<div class="region"><div class="contents">
<p class="p">To be able to disconnect someone who is viewing your desktop, you need to
 enable this option. If you select <span class="gui">Always</span>, this icon will be visible
 regardless of whether someone is viewing your desktop or not.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">If this option is disabled, it is possible for someone to connect to
 your desktop without your knowledge, depending on the security settings.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="sharing.html" title="Sharing">Sharing</a><span class="desc"> — 
      <span class="link"><a href="sharing-desktop.html" title="Share your desktop">Desktop sharing</a></span>,
      <span class="link"><a href="files-share.html" title="Dela ut och överför filer">Share files</a></span>…
    </span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
