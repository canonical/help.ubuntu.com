<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Kontakter</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Kontakter</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Använd <span class="app">Kontakter</span> för att spara, hantera eller redigera information om dina kontakter, lokalt eller i dina <span class="link"><a href="accounts.html.sv" title="Nätkonton">Nätkonton</a></span>.</p>
<div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="contacts-setup.html.sv" title="Starta Kontakter för första gången"><span class="title">Starta Kontakter för första gången</span><span class="linkdiv-dash"> — </span><span class="desc">Lagra dina kontakter i en lokal adressbok eller via ett nätkonto.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="contacts-connect.html.sv" title="Koppla ihop dig med din kontakt"><span class="title">Koppla ihop dig med din kontakt</span><span class="linkdiv-dash"> — </span><span class="desc">E-posta, chatta med eller ring en kontakt.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="contacts-add-remove.html.sv" title="Lägg till eller ta bort en kontakt"><span class="title">Lägg till eller ta bort en kontakt</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till eller ta bort en kontakt i den lokala adressboken.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="contacts-link-unlink.html.sv" title="Länka och avlänka kontakter"><span class="title">Länka och avlänka kontakter</span><span class="linkdiv-dash"> — </span><span class="desc">Kombinera information för en kontakt från flera källor.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="contacts-edit-details.html.sv" title="Redigera kontaktdetaljer"><span class="title">Redigera kontaktdetaljer</span><span class="linkdiv-dash"> — </span><span class="desc">Redigera informationen för varje kontakt.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="contacts-search.html.sv" title="Sök efter en kontakt"><span class="title">Sök efter en kontakt</span><span class="linkdiv-dash"> — </span><span class="desc">Sök efter en kontakt.</span></a></div>
</div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a><span class="desc"> — <span class="link"><a href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlöst</a></span>, <span class="link"><a href="net-wired.html.sv" title="Trådbundna nätverk">trådbundet</a></span>, <span class="link"><a href="net-problem.html.sv" title="Nätverksproblem">anslutningsproblem</a></span>, <span class="link"><a href="net-browser.html.sv" title="Webbläsare">webbsurfning</a></span>, <span class="link"><a href="net-email.html.sv" title="E-post &amp; e-postprogramvara">e-postkonton</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
