<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Nätverk, webb, e-post &amp; chatt</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Nätverk, webb, e-post &amp; chatt</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-grid ">
<div class="links-grid-link"><a href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="net-wireless-connect.html" title="Connect to a wireless network">Connect to wifi</a></span>,
      <span class="link"><a href="net-wireless-hidden.html" title="Connect to a hidden wireless network">Hidden networks</a></span>,
      <span class="link"><a href="net-wireless-edit-connection.html" title="Redigera en trådlös anslutning">Edit connection settings</a></span>,
      <span class="link"><a href="net-wireless-disconnecting.html" title="Why does my wireless network keep disconnecting?">Disconnecting</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-chat.html" title="Chatt &amp; sociala medier">Chatt &amp; sociala medier</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="net-chat-empathy.html" title="Snabbmeddelanden på Ubuntu">Chat on any network using <span class="app">Empathy</span></a></span>,
      <span class="link"><a href="net-chat-video.html" title="Video calls">make video calls</a></span>,
      <span class="link"><a href="net-chat-skype.html" title="Hur använder jag Skype på Ubuntu?">install skype</a></span>,
      <span class="link"><a href="net-chat-social.html" title="Social networking from the desktop">social networking apps</a></span>
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-mobile.html" title="Connect to mobile broadband">Connect to mobile broadband</a></div>
<div class="desc"><span class="desc">Connect to the internet using mobile broadband</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-email.html" title="E-post &amp; e-postmjukvara">E-post &amp; e-postmjukvara</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="net-default-email.html" title="Change which mail application is used to write emails">Default email apps</a></span>
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-security.html" title="Keeping safe on the internet">Keeping safe on the internet</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="net-antivirus.html" title="Behöver jag ett anti-virusprogram?">Antivirus software</a></span>,
      <span class="link"><a href="net-firewall-on-off.html" title="Enable or block firewall access">basic firewalls</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="contacts.html" title="Kontakter">Kontakter</a></div>
<div class="desc"><span class="desc">Kom åt dina kontakter.</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-general.html" title="Networking terms &amp; tips">Networking terms &amp; tips</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="net-findip.html" title="Hitta din IP-adress">Find your IP address</a></span>,
      <span class="link"><a href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?">WEP &amp; WPA security</a></span>,
      <span class="link"><a href="net-macaddress.html" title="What is a MAC address?">MAC addresses</a></span>,
      <span class="link"><a href="net-proxy.html" title="Define proxy settings">proxies</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-problem.html" title="Nätverksproblem">Nätverksproblem</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Troubleshooting wireless connections</a></span>,
      <span class="link"><a href="net-wireless-find.html" title="I can't see my wireless network in the list">finding your wifi network</a></span>…
        </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="sharing.html" title="Sharing">Sharing</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="sharing-desktop.html" title="Share your desktop">Desktop sharing</a></span>,
      <span class="link"><a href="files-share.html" title="Dela ut och överför filer">Share files</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-wired.html" title="Trådbunden anslutning">Trådbunden anslutning</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="net-wired-connect.html" title="Connect to a wired (Ethernet) network">Wired internet connections</a></span>,
      <span class="link"><a href="net-fixed-ip-address.html" title="Create a connection with a fixed IP address">Fixed IP addresses</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net-browser.html" title="Webbläsare">Webbläsare</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="net-default-browser.html" title="Change which web browser websites are opened in">Ändra förvald webbläsare</a></span>, <span class="link"><a href="net-install-flash.html" title="Install the Flash plug-in">installera Flash</a></span>, <span class="link"><a href="net-install-java-plugin.html" title="Install the Java browser plug-in">installera java-insticksprogrammet</a></span>, <span class="link"><a href="net-install-moonlight.html" title="Install the Silverlight plug-in">stöd för Silverlight</a></span>…</span></div>
</div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
