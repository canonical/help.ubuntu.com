<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns2="http://www.inkscape.org/namespaces/inkscape" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" height="500" id="svg10075" version="1.1" width="840" ns1:docname="gs-goa2.svg" ns2:version="0.92.4 5da689c313, 2019-01-14">
  <ns0:defs id="defs10077">
    <ns0:linearGradient id="RHEL7" ns3:paint="gradient">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop id="stop11074" offset="0" style="stop-color:#eeedec;stop-opacity:1;"/>
      <ns0:stop id="stop11076" offset="1" style="stop-color:#eeedec;stop-opacity:1"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop id="stop7012" offset="0" style="stop-color:#eeedec;stop-opacity:0;"/>
      <ns0:stop id="stop7014" offset="1" style="stop-color:#eeedec;stop-opacity:0"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" gradientUnits="userSpaceOnUse" id="linearGradient7064" x1="-18.33782" x2="713.42853" y1="490.54935" y2="490.54935" ns2:collect="always" ns4:href="#GNOME"/>
    <ns0:filter color-interpolation-filters="sRGB" height="1.1308649" id="filter5601" width="1.2058235" x="-0.10291173" y="-0.065432459" ns2:collect="always">
      <ns0:feGaussianBlur id="feGaussianBlur5603" stdDeviation="0.610872" ns2:collect="always"/>
    </ns0:filter>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient5885" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns2:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop id="stop5718" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17441" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns2:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop id="stop17445" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop17447" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17453" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns2:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17455" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns2:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient ns2:collect="always" ns4:href="#linearGradient5716" id="linearGradient1244" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient ns2:collect="always" ns4:href="#linearGradient5716" id="linearGradient1246" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
  </ns0:defs>
  <ns1:namedview bordercolor="#666666" borderlayer="true" borderopacity="1.0" fit-margin-bottom="0" fit-margin-left="0" fit-margin-right="0" fit-margin-top="0" height="0px" id="base" pagecolor="#eeeeec" showgrid="false" width="0px" ns2:current-layer="g6301" ns2:cx="24.172052" ns2:cy="234.91841" ns2:document-units="px" ns2:pageopacity="1" ns2:pageshadow="2" ns2:showpageshadow="false" ns2:window-height="1403" ns2:window-maximized="1" ns2:window-width="2560" ns2:window-x="3440" ns2:window-y="0" ns2:zoom="1" ns2:document-rotation="0">
    <ns2:grid empspacing="5" enabled="true" id="grid17504" snapvisiblegridlinesonly="true" type="xygrid" visible="true"/>
  </ns1:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g id="layer1" transform="translate(0,-992.3622)" ns1:insensitive="true" ns2:groupmode="layer" ns2:label="bg">
    <ns0:rect height="656" id="background" style="fill:url(#BLANK);" width="866" x="-16" y="855.36218" ns2:label="background"/>
  </ns0:g>
  <ns0:g id="layer2" transform="translate(0,-540)" ns2:groupmode="layer" ns2:label="fg">
    <ns0:g id="g11020" transform="translate(-81,-139.36217)">
      <ns0:circle id="path11014" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;enable-background:accumulate" transform="translate(2,453.36217)" cx="120" cy="278" r="17"/>
      <ns0:text id="text11016" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" xml:space="preserve"><ns0:tspan id="tspan11018" x="122.29289" y="736.36218" ns1:role="line" style="font-size:14px;line-height:1.25">3</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:path ns2:connector-curvature="0" ns1:nodetypes="sssccccss" style="fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:5.36666679;stroke-miterlimit:4;stroke-opacity:1" id="path5430" d="m 141.41664,1245.6834 h 561.16668 c 5.94626,0 10.73333,4.8289 10.73333,10.8272 v 329.4895 H 702.58332 141.41664 130.68331 v -329.4895 c 0,-5.9983 4.78707,-10.8272 10.73333,-10.8272 z"/>
    <ns0:path ns2:connector-curvature="0" style="fill:none;stroke:#000000;stroke-width:2.72237611;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" id="path5361" d="m 132.16207,1295.6167 c 570.10453,0 580.39987,0 580.39987,0"/>
    <ns0:g transform="matrix(1.262736,0,0,1.262736,678.32655,1261.9854)" style="fill:#0c0000;fill-opacity:1" id="g5363">
      <ns0:g transform="translate(-60,-518)" style="display:inline;fill:#0c0000;fill-opacity:1" id="g5365"/>
      <ns0:g transform="translate(-60,-518)" style="fill:#0c0000;fill-opacity:1" id="g5367"/>
      <ns0:g transform="translate(-60,-518)" style="fill:#0c0000;fill-opacity:1" id="g5369"/>
      <ns0:g transform="translate(-60,-518)" style="fill:#0c0000;fill-opacity:1" id="g5371">
        <ns0:g transform="translate(19,-242)" style="display:inline;fill:#0c0000;fill-opacity:1" id="g5373">
          <ns0:path ns2:connector-curvature="0" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.78124988;marker:none;enable-background:new" id="path5375" d="m 45,764 h 1 c 0.01037,-1.2e-4 0.02079,-4.6e-4 0.03125,0 0.254951,0.0112 0.50987,0.12858 0.6875,0.3125 L 49,766.59375 51.3125,764.3125 C 51.578125,764.082 51.759172,764.007 52,764 h 1 v 1 c 0,0.28647 -0.03434,0.55065 -0.25,0.75 l -2.28125,2.28125 2.25,2.25 C 52.906938,770.46942 52.999992,770.7347 53,771 v 1 h -1 c -0.265301,-10e-6 -0.530586,-0.0931 -0.71875,-0.28125 L 49,769.4375 46.71875,771.71875 C 46.530586,771.90694 46.26529,772 46,772 h -1 v -1 c -3e-6,-0.26529 0.09306,-0.53058 0.28125,-0.71875 l 2.28125,-2.25 L 45.28125,765.75 C 45.070508,765.55537 44.97809,765.28075 45,765 Z"/>
        </ns0:g>
      </ns0:g>
      <ns0:g transform="translate(-60,-518)" style="fill:#0c0000;fill-opacity:1" id="g5377"/>
      <ns0:g transform="translate(-60,-518)" style="fill:#0c0000;fill-opacity:1" id="g5379"/>
      <ns0:g transform="translate(-60,-518)" style="fill:#0c0000;fill-opacity:1" id="g5381"/>
    </ns0:g>
    <ns0:text xml:space="preserve" y="1274.9995" x="427.99988" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:32.20000076px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2.6833334" id="text12012"><ns0:tspan style="font-size:13.99999905px;line-height:1.25;stroke-width:2.6833334" ns1:role="line" y="1274.9995" x="427.99988" id="tspan12014">Nätkonton</ns0:tspan></ns0:text>
    <ns0:rect y="1416.7651" x="189.79674" height="169.23441" width="484.75693" id="rect884" style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1"/>
    <ns0:g ns2:label="#g5607" transform="matrix(2.7589319,0,0,2.7589319,485.15811,1476.7641)" style="display:inline" id="default-pointer-c">
      <ns0:path ns2:connector-curvature="0" ns1:nodetypes="cccccccc" style="color:#000000;display:block;overflow:visible;visibility:visible;opacity:0.6;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;filter:url(#filter5601);enable-background:accumulate" id="path5567" d="M 27.135224,2.8483222 V 19.288556 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z"/>
      <ns0:path ns2:connector-curvature="0" ns1:nodetypes="cccccccc" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17453);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" id="path5565" d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z"/>
      <ns0:path ns2:connector-curvature="0" ns1:nodetypes="cccccccc" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17455);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" id="path6242" d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z"/>
    </ns0:g>
    <ns0:g ns2:label="go-previous" transform="translate(46.922014,743.97752)" style="display:inline" id="g4705">
      <ns0:rect y="518" x="-116" width="16" transform="scale(-1,1)" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none;enable-background:new" id="rect10837-5-8-1" height="16"/>
      <ns0:path ns2:connector-curvature="0" ns1:nodetypes="ccsccccccccccc" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.78124988;marker:none;enable-background:new" id="path10839-9-9-5" d="m 112.01352,520 h -1 c -0.0104,-1.2e-4 -0.0208,-4.6e-4 -0.0313,0 -0.25495,0.0112 -0.50987,0.12858 -0.6875,0.3125 l -6.29767,5.71875 6.29772,5.71875 c 0.18816,0.18819 0.45346,0.28125 0.71875,0.28125 h 1 v -1 c 0,-0.26529 -0.0931,-0.53058 -0.28125,-0.71875 l -4.82897,-4.28125 4.82897,-4.28125 c 0.21074,-0.19463 0.30316,-0.46925 0.28125,-0.75 z"/>
    </ns0:g>
    <ns0:rect y="1254.469" x="139.53026" width="31.999998" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.99999994;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" ry="3.9999998" rx="3.9999998" id="rect15386" height="31.999998"/>
    <ns0:rect ry="3.5355337" rx="3.5355337" y="1306.4878" x="696.37891" height="121.62237" width="7.0710673" id="rect977" style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal"/>
    <ns0:rect style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1" id="rect979" width="40.955532" height="39.882473" x="214.06105" y="1437.2712"/>
    <ns0:rect y="1497.2714" x="214.06105" height="39.882473" width="40.955532" id="rect981" style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1"/>
    <ns0:rect style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1" id="rect983" width="40.955532" height="28.728062" x="214.06105" y="1557.2715"/>
    <ns0:rect y="1446.675" x="270.11478" height="19.79899" width="178.1909" id="rect985" style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal"/>
    <ns0:rect style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect987" width="127.27921" height="19.79899" x="270.11478" y="1505.3649"/>
    <ns0:rect y="1565.469" x="270.11478" height="14.469899" width="203.64674" id="rect989" style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal"/>
    <ns0:flowRoot style="font-style:normal;font-weight:normal;font-size:40px;line-height:1.25;font-family:sans-serif;letter-spacing:0px;word-spacing:0px;fill:#000000;fill-opacity:1;stroke:none" id="flowRoot1005" xml:space="preserve" transform="matrix(2.6833333,0,0,2.6833333,-1275.5101,-1072.8539)"><ns0:flowRegion id="flowRegion1007"><ns0:rect y="199" x="186" height="122" width="488" id="rect1009"/></ns0:flowRegion><ns0:flowPara id="flowPara1011"/></ns0:flowRoot>    <ns0:text id="text1074" y="1403.0002" x="192.0002" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:14.66666794px;line-height:1.25;font-family:sans-serif;-inkscape-font-specification:'sans-serif, Normal';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.99999994" xml:space="preserve"><ns0:tspan style="stroke-width:0.99999994" y="1403.0002" x="192.0002" id="tspan1072" ns1:role="line">Lägg till ett konto</ns0:tspan></ns0:text>
    <ns0:g ns2:label="account-facebook" transform="matrix(2.5,0,0,2.5,-155.93914,436.27124)" style="display:inline;stroke-width:0.80000001" id="g3922">
      <ns0:rect ns2:label="audio-volume-high" y="20" x="-194" width="16" transform="rotate(-90)" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.80000001;marker:none" id="rect2941" height="16"/>
      <ns0:path ns2:connector-curvature="0" ns1:nodetypes="sssscccccscccsscccccsssss" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.40000001;marker:none;enable-background:new" id="rect14063" d="M 22.116732,178 C 20.946094,178 20,178.94979 20,180.125 v 11.75 c 0,1.17521 0.946094,2.125 2.116732,2.125 h 6.910506 v -6 h -0.99611 v -2 h 0.99611 v -1.0625 c 0,-1.84445 1.374066,-2.88912 3.175096,-2.9375 h 1.77432 v 2 H 32.88716 c -0.625856,0 -0.902724,0.22291 -0.902724,0.90625 V 186 h 1.712062 l -0.217898,2 h -1.494164 v 6 h 1.898832 C 35.053906,194 36,193.05021 36,191.875 v -11.75 C 36,178.94979 35.053906,178 33.883268,178 Z"/>
    </ns0:g>
    <ns0:path ns2:connector-curvature="0" ns1:nodetypes="ccccscscccccscccsccssscccccsccccsccccccccsccc" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.49999997;marker:none;enable-background:new" id="path14750" d="m -94.36077,823.29363 -4.452965,-0.0161 c -3.138825,1.63525 -3.608415,5.71553 -2.578065,9.45277 1.36187,4.93932 4.083657,8.40395 7.734144,7.26542 5.092108,-1.58856 5.241113,-5.74711 3.671739,-10.62463 -0.830009,-2.57976 -2.369518,-4.65822 -4.374853,-6.07402 z m 12.421472,7.71456 c 0,2.19931 -0.894865,4.07649 -1.874926,5.54669 v 0.0786 l -0.234523,0.15617 c 0,0 -0.636862,0.74801 -1.406201,1.48437 -0.768238,0.73649 -1.953064,1.7187 -1.953064,1.7187 -0.964095,0.72458 -1.484286,1.68245 -1.484286,2.73423 0,1.05541 0.670619,2.00936 1.640563,2.73429 0,0 1.966911,1.20517 3.046764,2.10935 1.079398,0.90471 2.343704,2.10928 2.343704,2.10928 1.461961,1.37465 2.421762,3.56524 2.421762,6.01542 0,2.1102 -0.669116,4.02371 -1.796814,5.39044 l -1.718701,2.18745 h 10.702743 c 2.926551,0 5.312356,-2.37442 5.312356,-5.31235 v -29.37402 c 0,-2.9379 -2.385805,-5.3123 -5.312356,-5.3123 -1.434564,-0.0134 -4.553536,0.003 -4.553536,0.003 l -0.03837,2.464 -6.414723,0.71948 c 0.93863,1.63007 1.295782,3.25706 1.319878,4.5464 z m -24.999192,6.09358 v 14.06201 c 4.34099,-2.90643 12.108995,-2.96866 12.108995,-2.96866 0,0 0.03354,-0.0469 0,-0.0786 -3.114384,-2.39415 -1.796813,-5.15624 -1.796813,-5.15624 -4.815402,0.41026 -7.016572,-1.38709 -10.312182,-5.85914 z m 12.655885,13.82767 c -4.326311,0.24311 -9.893045,2.03421 -9.999685,6.32789 0,2.56833 1.67199,4.89633 4.06233,5.93731 0,0 0.0859,0.055 0.15617,0.0786 h 0.07862 11.327745 c 0,0 0.02147,-0.1119 0.07862,-0.15617 6.127821,-5.42329 1.500386,-8.5677 -3.749905,-12.10895 -0.09526,-0.0633 -0.234523,-0.0786 -0.234523,-0.0786 -0.54748,-0.0215 -1.100676,-0.0344 -1.718675,0 z"/>
    <ns0:path style="display:inline;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:5.36666679;stroke-miterlimit:4;stroke-opacity:1" d="M 83.416662,568.68327 H 776.58334 c 5.9463,0 10.73334,4.78707 10.73334,10.73333 v 432.6333 H 776.58334 83.416662 72.683329 V 579.4166 c 0,-5.94626 4.787067,-10.73333 10.733333,-10.73333 z" id="path5430-2" ns2:connector-curvature="0" ns1:nodetypes="sssccccss"/>
    <ns0:path ns2:connector-curvature="0" id="path5361-7" d="M 74.162087,618.61661 H 786.56199" style="display:inline;fill:none;stroke:#000000;stroke-width:2.72237611;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns1:nodetypes="cc"/>
    <ns0:path style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3.58466077;marker:none;enable-background:new" id="path5375-0" d="m 754.37986,585.03757 h 2.01245 c 0.0215,-2.4e-4 0.0419,-9.4e-4 0.0628,0 0.51308,0.0215 1.02608,0.25867 1.38355,0.62889 l 4.59089,4.59086 4.65376,-4.59086 c 0.53454,-0.46387 0.89891,-0.6148 1.38355,-0.62889 h 2.01245 v 2.01245 c 0,0.57648 -0.0692,1.10813 -0.50313,1.50932 l -4.59086,4.59088 4.52799,4.528 c 0.3787,0.37867 0.56597,0.91254 0.566,1.44645 v 2.01242 h -2.01245 c -0.5339,0 -1.06778,-0.1873 -1.44645,-0.566 l -4.59086,-4.59089 -4.59089,4.59089 c -0.37867,0.37873 -0.91257,0.566 -1.44645,0.566 h -2.01245 v -2.01242 c 0,-0.53391 0.1873,-1.06778 0.56603,-1.44645 l 4.59086,-4.528 -4.59086,-4.59088 c -0.42413,-0.39169 -0.61011,-0.94435 -0.56603,-1.50932 z" ns2:connector-curvature="0" ns1:nodetypes="ccccccccscccccscccscsccccc"/>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:32.20000076px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2.6833334" x="519.99988" y="597.99994" id="text12012-9"><ns0:tspan ns1:role="line" id="tspan12014-3" x="519.99988" y="597.99994" style="font-size:13.99999905px;line-height:1.25;stroke-width:2.6833334">Nätkonton</ns0:tspan></ns0:text>
    <ns0:g id="g9286" transform="matrix(2.6833333,0,0,2.6833333,-1322.5101,-1214.8539)">
      <ns0:g id="g3921" transform="matrix(0.37267081,0,0,0.37267081,493.07637,552.48134)" style="display:inline"/>
    </ns0:g>
    <ns0:rect width="15.999999" height="15.999999" x="-103.92204" y="584.97754" id="rect10837-5-8-1-6" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.99999994;marker:none;enable-background:new" transform="scale(-1,1)"/>
    <ns0:path d="m 99.935584,586.97746 h -0.999998 c -0.01073,-1.1e-4 -0.02147,-4.6e-4 -0.0314,0 -0.254917,0.0107 -0.50986,0.12853 -0.687497,0.3125 l -6.297676,5.71875 6.29773,5.71874 c 0.188102,0.1881 0.453456,0.28127 0.718758,0.28127 h 0.999997 v -1 c 0,-0.26538 -0.09311,-0.5306 -0.28124,-0.71876 l -4.82898,-4.28125 4.82898,-4.28124 c 0.210642,-0.19454 0.303136,-0.46926 0.28124,-0.75001 z" ns2:connector-curvature="0" id="path10839-9-9-5-0" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.78124988;marker:none;enable-background:new" ns1:nodetypes="ccsccccccccccc"/>
    <ns0:rect style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.99999994;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" id="rect15386-6" width="31.999998" height="31.999998" x="80.530251" y="577.46942" rx="3.9999998" ry="3.9999998"/>
    <ns0:text id="text946" y="597.99994" x="177.99998" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:32.20000076px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2.6833334" xml:space="preserve"><ns0:tspan style="font-size:13.99999905px;line-height:1.25;stroke-width:2.6833334" y="597.99994" x="177.99998" id="tspan944" ns1:role="line">Inställningar</ns0:tspan></ns0:text>
    <ns0:rect transform="scale(-1,1)" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.99999994;marker:none;enable-background:new" id="rect948" y="584.97754" x="-268.92215" height="15.999999" width="15.999999"/>
    <ns0:rect ry="3.9999998" rx="3.9999998" y="577.46942" x="245.53044" height="31.999998" width="31.999998" id="rect952" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.99999994;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate"/>
    <ns0:g ns2:label="open-menu" id="g7352" transform="translate(233.9223,309.97744)" style="display:inline;enable-background:new">
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" id="rect7354" width="16" height="16" x="20" y="276"/>
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7356" width="9.9996014" height="2.0002136" x="23.000198" y="278.99979"/>
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7358" width="9.9996014" height="2.0002136" x="23.000198" y="282.99979"/>
      <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7360" width="9.9996014" height="2.0002136" x="23.000198" y="286.99979"/>
    </ns0:g>
    <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:15.99999905;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7822" width="212.00002" height="45.999996" x="73.999947" y="661"/>
    <ns0:text id="text7826" y="687.99988" x="125.57443" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:32.20000076px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2.6833334" xml:space="preserve"><ns0:tspan style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:13.99999905px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;text-anchor:start;fill:#ffffff;stroke-width:2.6833334" y="687.99988" x="125.57443" id="tspan7824" ns1:role="line">Nätkonton</ns0:tspan></ns0:text>
    <ns0:path style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" d="M 286.53042,567.46946 V 1010" id="path7828" ns2:connector-curvature="0"/>
    <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7830" width="48" height="9" x="125.00006" y="636"/>
    <ns0:rect y="725.99994" x="125.00006" height="9" width="48" id="rect7832" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
    <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7834" width="48" height="9" x="125.00006" y="766"/>
    <ns0:rect y="766" x="185.00018" height="9" width="77" id="rect7836" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
    <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="path7840" cx="97.581062" cy="641.03552" r="11.418957"/>
    <ns0:circle r="11.418957" cy="732.03546" cx="97.581062" id="circle7842" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
    <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.99999994;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle7844" cx="97.581062" cy="770.03546" r="11.418957"/>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:21.33333397px;line-height:1.25;font-family:sans-serif;-inkscape-font-specification:'sans-serif, Normal';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1" x="420" y="1351" id="text1050"><ns0:tspan ns1:role="line" id="tspan1048" x="420" y="1351">Anslut till dina data i molnet</ns0:tspan></ns0:text>
    <ns0:rect style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1" id="rect1212" width="450.75693" height="268.23441" x="309.55975" y="741.81555"/>
    <ns0:g id="g1220" style="display:inline" transform="matrix(2.7589319,0,0,2.7589319,597.92114,801.81449)" ns2:label="#g5607">
      <ns0:path d="M 27.135224,2.8483222 V 19.288556 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path1214" style="color:#000000;display:block;overflow:visible;visibility:visible;opacity:0.6;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;filter:url(#filter5601);enable-background:accumulate" ns1:nodetypes="cccccccc" ns2:connector-curvature="0"/>
      <ns0:path d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path1216" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient1244);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" ns1:nodetypes="cccccccc" ns2:connector-curvature="0"/>
      <ns0:path d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path1218" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient1246);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" ns1:nodetypes="cccccccc" ns2:connector-curvature="0"/>
    </ns0:g>
    <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect1222" width="7.0710673" height="121.62237" x="771.49097" y="628.61664" rx="3.5355337" ry="3.5355337"/>
    <ns0:rect y="882.32166" x="326.82407" height="39.882473" width="40.955532" id="rect1224" style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1"/>
    <ns0:rect style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1" id="rect1226" width="40.955532" height="39.882473" x="326.82407" y="942.32178"/>
    <ns0:rect y="1002.3219" x="326.82407" height="9.7280617" width="40.955532" id="rect1228" style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1"/>
    <ns0:rect style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect1230" width="178.1909" height="19.79899" x="382.87781" y="891.72546"/>
    <ns0:rect y="950.41528" x="382.87781" height="19.79899" width="127.27921" id="rect1232" style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal"/>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:14.66666794px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.99999994;" x="311.76321" y="728.05066" id="text1238"><ns0:tspan ns1:role="line" id="tspan1236" x="311.76321" y="728.05066" style="stroke-width:0.99999994;-inkscape-font-specification:Cantarell;font-family:Cantarell;font-weight:normal;font-style:normal;font-stretch:normal;font-variant:normal;">Lägg till ett konto</ns0:tspan></ns0:text>
    <ns0:text id="text1242" y="676.05042" x="532.763" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:21.33333397px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1" xml:space="preserve"><ns0:tspan y="676.05042" x="532.763" id="tspan1240" ns1:role="line">Anslut till dina data i molnet</ns0:tspan></ns0:text>
    <ns0:rect style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1" id="rect1248" width="40.955532" height="39.882473" x="326.82407" y="762.43909"/>
    <ns0:rect y="822.43921" x="326.82407" height="39.882473" width="40.955532" id="rect1250" style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:1;stroke-opacity:1"/>
    <ns0:rect y="771.8429" x="382.87781" height="19.79899" width="178.1909" id="rect1252" style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal"/>
    <ns0:rect style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:20;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect1254" width="127.27921" height="19.79899" x="382.87781" y="830.53271"/>
    <ns0:g transform="translate(-120.9999,206)" id="g6301" ns2:label="goa-panel" style="enable-background:new">
      <ns0:path style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.99999976;marker:none;enable-background:accumulate" d="M 101 137 A 4.0000017 4.0000017 0 0 0 97.369141 139.33398 A 2.9999998 2.9999998 0 0 0 96 139 A 2.9999998 2.9999998 0 0 0 93 142 A 2.9999998 2.9999998 0 0 0 93.181641 143.02344 A 2.5 2.5 0 0 0 91 145.5 A 2.5 2.5 0 0 0 93.5 148 L 104 148 A 3.0000013 3.0000013 0 0 0 107 145 A 3.0000013 3.0000013 0 0 0 104.83594 142.12109 A 4.0000017 4.0000017 0 0 0 105 141 A 4.0000017 4.0000017 0 0 0 101 137 z " transform="translate(120.9999,334)" id="circle3296"/>
      <ns0:rect width="16" height="16" x="211.9998" y="468" id="rect3664" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1.78100002;marker:none;enable-background:new"/>
    </ns0:g>
  </ns0:g>
</ns0:svg>
