�PNG

   IHDR     }   `��  �zTXtRaw profile type exif  xڭ�ir9F��sl�Hk��`�?/���-��c{H���UXr��R8�����QzΡJ3�G������x^S��������?�~_�9Tx/�?M�~_�m��'��@��_����=�}�=Q�e>��{��__�� 㵭���߷0���c#O��2?����O�F��0O���T"�������P:�����?F����
�Wq�����R�'}��o�>e�}�s�j~�R>Y��y<$�:+O��6s�����q>�׊>E���v�=��Q�P�{S[|>q�d$��K����hϳ�4�zQ
;�8y��S&]7մ�H7��}��k>!7>�ryZi��E&ɢ?�͍��b�s=i�%[Kz��q�g6c�85'KO��3���z+��l���.����@�WN##龃*O�?����B�ģ�-�	�|1%���It�D��Ճ	�x@��ZXL*d���"ISl9�������3=3�@ɛE�Z���>5�����%s8p0#R�4rCߑ�Z��iը�!E���41�2�hUQզ���VC���5k�+VML��Y��s/��t�[�}��<�zp�3�2�0u�i�ϱ(�U�,]m��k��?��m�=N:�ҩG��v��3.�vK����ۮ�~Ƿ���������Y�O����-km�c��p"�3�$2�<t��EK�fϜ�,�LWHf��9��3F�IYn��]ȯ�z��(o����7s�S����1o_em;�'c�.���B�ݼ���t�M���C��2v_gɹ�)qUm�\*����\ �X�'����¸(n�+y�Z��}�k�0���w��8���������tuT��9[���OQ;b��V5˃����Mg�o�����;�t�r�v5@��=3�7�yr���kj�X֦�h?��D͔�ړ+����K_Ųٺj�:ݾ�i7݇�B�g��S
��4�������PI*�=˱F Xm��u 6�ᔪs�9��r��Y+��QVki�fFt�(�M�n��N`��4�����	Qf�;��M�X��.Y�ZZ��Ѿ�g*�P3��r���b�"ZV�L�jПH�J=�ZL�ã&
�,�YX>���X,��ni�Ǌ�GBtZas�Ls��r3�|�N��DEg���4��Yr�3�mD���d�3{pA�m��g��N(Cj���Z�bzYS�m�!�k?*L��]�7� w�3�$�<�en�K�X{�+K��Tg1��48Y�ܐ��űZH�������n>i殥P�Q�hf`˶a%^�Q�~� �
ᴵFkz�>8�`_�Cq������/	��i`�h_��w�BY���]�|��E�c�|d��ѷV�|ս��I[����-qf�M�{:�e[�i��p�\�N�6]��i�L���^�����^=0�`=������o���|A8@.@V��XD4
�����-����^*���֏�ej ����Δ�A����E�*�W�8�I>qoY��;l�
�k��>�Rҗ�EU�!Ӿ����T���Pn����h85����~Ԋ������\R.��^��;;�D1��{=g�Y�e��� ���~f��`��|s�z�:8.�@z�~�B1�B��/��U)�P�ke���ܧl9�|:JQ�S�2�u�t�9�c.y�E�xD'1�^0+pE���R�3��X��	�����
-�:*}0Aaѵ�-C���&Z��S[g�,��D�%�`Ђ��z7Ox<A���@����0)���xU�FC0ą+(�����iAE�z�d��������h�2w����MKr99R����g��C��މYvJ�%�@��ҋ�"��9���K��ں˳J`1
�$��R�=�@��ᣏ��@��2��}�A�{�-+\��;�I8�>�w���[�n�ꃿ�Â/�#��LM�
��9�Ƹ�ѓ|�X�J��^����h�HY6H�%��u����,ә#���f�!��N�־�A�9!>/־(��t�V8�vc,G��.�́%�a@B�긃�R�(�z Aݫ��rd"���6 �?�M�i�do��v��̣^��W�^�Y`F��D�n��t�8"j�XA�tQ ��T$g)��@N8!ĎB���k�#��g 3QS�а�ʞl T������'��y�M�7F���s������9�C)��IL3�U�����XB�`VsQ�ܷ�rΫ���j���� ׽ q���9ھ���u�}aA���V���������G{��+d8����Ӟ����>#�]��?9񋍼�v��j�����v�W���톟M��v%_�������<+� B�����h �0 �;y������l8���F�	/Ӱ�t��O�%�fA���:Z����X���Ԅ_YoO�2c�I�PԆN
zr�5'	�N�@o�ʺ�u!rB�%
����E�3���a�p����^�A���m�����.�D��U��>��������f���l�8�C@�D4�5�&"����(�w\�8�c�15{��٬�3|춌��h�Ӱ�!rn�˨�z}ga�0�r�ࡋ�bȝ)���A�АK�`� �9���~0��j@������8��4p� 6�]�sG=t�J�p���&V1��)c˰2��i����@���t��(>�ZW��# h�El@��|�|K9�(W*��%c��V���J�@V��s&5���|7��D�ķ�auq��[!��+V�%����_9���� �uF��1�{�]�´C��..�؇�r\�4��|���No8�-{p�'5�����2��.A�.�jb����C��Acj��,tg�rt^#J��	�cرN]
[Į��3�� ������#�	q�J6�w7E�.�=W(Ń+�D}*dd(��}�݅�vռP�Q��>�Ơ�����-~w��|�m� �}+�
 ��$�4�����0���v��ˎ87�g�+�N.m�\P�ب3:7��*���!8��,8A
q,�����>2JVx��d���ל=�d����`��b(r��8V%f��$�
�z@1��C�c���{�:9��������э�c���5խ#�E��F�k�T�^�ܜeO��?���ރV"���i~1��|����=�(d�	�=���#�j[J�Κ�˰����K��\�����;LxNE�x���܇FH>)Fɹ�2'�2���:P셁A���8� �����<j낌��7���_R�:�.\�(�Q�?k*���-Dack-����Ub|\`@)�M�{D���E����4B�G�u��d��C��;�.���N�Ro���.�~<m�{�`@F2�!of��x����`�G�>��������O�������2�;�����Wï��`4�fd�O��24�zVT��b<Z�{� L��֟I��/���?��|�{�������!�I  �iCCPICC profile  x�}�=H�@�_S�*U3�8D�NDE�
E�j�V�G��IC���(��X�:�8���*� �NN�.R���B����������J�f���n��xLHgV��+����˘�|��=l���,�s�5k)@@ �U�&� �޴��ļR�T�s�1�.H��t��7�y�9�ɛ��<1O,�[Xna�`j�S�U�)�K{�2�b��*J��ᬾ��t�C�cK!@FE�`#J�N��$��|���_$�L�"r,�������Z��	/)�_�c����|;N�>Wz�_�3��W�Z���.����\� O�dJ����r��}S��׼��8} R�U�88F��������=���<er�ԏ��  xiTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:85010c16-09b1-4807-aab2-f1ebfb4c8b30"
   xmpMM:InstanceID="xmp.iid:11e864dc-a74a-4b71-9f67-6c3aec0f2647"
   xmpMM:OriginalDocumentID="xmp.did:5fdf32e5-48b9-4b9e-8ce3-6ea3aa5ab3cc"
   dc:Format="image/png"
   GIMP:API="2.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1663187632836218"
   GIMP:Version="2.10.32"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP 2.10"
   xmp:MetadataDate="2022:09:14T22:33:52+02:00"
   xmp:ModifyDate="2022:09:14T22:33:52+02:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:ceed33a4-9b2a-4a76-84fd-c0555202e9fe"
      stEvt:softwareAgent="Gimp 2.10 (Linux)"
      stEvt:when="2022-09-14T22:33:52+02:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>�3-   bKGD � � �����   	pHYs  �  ��+   tIME�
!�2I  IDATx��{Tg���L.���N$��T.QQ.��Pѵ��s���U����gm�Z�u{j�=kʶ���h�k=���T�`Q�V�6�Z/�EA	$\�2���i
��h��_��w�ɼy�y/���aEFF"  �  @K  Z �  �% x�p��=��j6����n�Xz�'[�V��⭷�Z�xqHH�ٳg�O;n�8�Hd0��=�\������ŋ�?���.EGGGFFr8N�x��3f�t:(Y �� ���H����E%''wtt���uvv���(�J����WBBB�̙3.������Dooo��|�������������k׮9�N�T���kjjp�����x������F??�ѣG{yyq�\�����߻��gRK���F�����cccI�DUWW����6l�"���C%$$DFF~��b��k�X��׿�>}ڝω'���I������v�k��v�ڵ ��ZmAA��Z�`Acc�G}4f��װZ�+V��r�
���S�C������ر�O>A'&&n߾��K�.�_�~���\.���>��_|�Ezzz^^EQ[�l�D�|�L�r�ر��/_>p����
ǚ�={6�źr�ʵk�BEEE˖-�9s�ܹsO�:%�V�Z���k�믿��/������qRVV���Bw��9t�СC�ƍGQB�d2M�6��t"��R�q���?~�o�ۮ]�JKK�޽���9s� �222�DNy��ш��?�����ٸ3����0�o��v�]"�p���i�R)�x�7<�c%`*++=&%%͚5���4  �f�9r����O�T���|9,T x���0L����!��_cc#N�����ԄwR�����7'N�hnn���Y�nB�ȑ#V�!4q�D�R���5g��ñj�*��g^K}R__�JJJھ}�^�ߺukMMMPPп�����B����:m�4O9y�r�:�|��c�zv����B</;;���mѢE���d��'{��9s�M�S�NMLLt�\�ӟ���CBB�y睷�z+==]�����ؿ?n����.]��w�>}�����%K�̝;׭1 xz`=�w�\������4�=:u�B�PP���@�4�r��% �>  �%  - h	 @K  ��  � �%  @K  Z������������f�Z��b�D"�T�����Ҁ`�h4Z,�J��j�K�V���������(�J�b����ă��BHw��!"**J�T��|� ����r�����h4������A���ˋ �����M?��U�.���[j�h4A}��P�����6���Dœ����7vvv��չw���D"l�����ɱc�.\�����f��b����1�n�X�װ,\�0**jɒ%���w��u��)��S:^jkkS�Tl6�OC�_ZC6���'�qH,������|��#F�p����$���F����q��Y��įn��INN�h4V��ҥK7o�D�L&l&�	���oii���o=��h4			\.��~�'"��������B�ĉ+**���v�j���rz (�>]f͚���KKKϟ?��K/=�����?���?Θ1���111�{��w�~��W5M\\��ￏ��Y�f�̙x{�����틎�NII���w�N������###��ݻp�B�?'''77��?����j}��������o�0|>�O�y��!����V�^������������lٲ���+Vx&3f������|�	6��v���۷�޽!�h�"�;�f�׭[WPP����*//���-))1�L!oo����;�C�ci�B̀�}�Q���ÿ��k�Pii)EQ�&M��r4M����^���wߍ��	

�=b��sss'O�L�d�����k4��⏇�~~~�f����cqq1�0�W��=
Bc���p�����f��v��7o��j]�l����1o޼�g>��S>�_\\\UU8a	��ۗ.]�hѢ��\�L��_n߾�3�bZ���b���r�ݳ�����
��� ��ՒP(4�LB���){'�p8���f��)++��̔J��
��F3q����d\�333�Lv���6 �&L����������~r���Ah�چ�����/��F��2������B�@�R�D9���xR��d29���{wN��d2I$�s�N�*
�{�O�y�f�ٌ�����p03j�(��J�Z�ti�z��w�ܡi��8�`0�t���,�L9++�ojj:w�\vv6v����6�Z
xB�I�E�����xRWWGQ9�f�ܹǏ���f�ȑ#/��Ҟ={�̧��e�Ν��������������J�'�|B�tkk�J���Ϫ��z�ٴiS^^^YYM���lxnn�m���˝N��n��q�0�z<���l����h���ݷoߦiZ����0��C�B���p?GX�؂$I��`���f�ȑf���@H��p8����B.�����b���r�D"�dC{{��l�(J�T�1	 �� �0�����f�����
�DB�$,`�4`��X|>����*@K�(� � h	 @K  Z  � �%  - h	  � <y� �b-�2���x �ڇ�"�@�b�p��ۃ:�E�\���1���xtdubb����i�1g�#�V�e���{���q�\�P�=�{��+��b��s�4Fzt�ѣ�x{{GFF䊱�1~~�'_p���w�4@�x��=�y<^@���ǏO�6M"����<�r�j��d2��|�'�����\.�^����imms6h�����$�#��\^s����8���������.��h�6Iv���x�\��j:;m�n���p9l_�T�pt���Vk'T8h�ʣ{ ��[,���:�^��@%###((�n���j�@�����2e����;qjj�B!G�T�^V(�3f̘0a� ��b͙3;&�����N�:�0aB@@ �9o�K���#G�HOOw����!��~��������A�4P�944�ݸQ5~��.x�&����Ҫ��~��G��իWCB�kkk/_~�;~RRbEEeee%BH$�͟?���j�f�?R�T�T�ڵ�~sA��ǟ;w�ҥK������?������)::*66��o�@��vi�<��B!W*�UU7Buuu<W��e,�V{gd���tXHG,�p3������P(�V����@ε�l.�+))��Ϗ�a������7n��7nTyEPP���q			j�Z&�C��vi��=�rhh��錎�r�d���b;U��R�Dݽ{w��J$�B��~n�67���T��p8�:"blRR"I��/_9�|�Ÿ���KOO�p8��5&�Y&�j4�p����Z�C{ |�v���s��u�VXXI������U�;{v�7�q�$3��/ϩ�N'��qOc`�>�_y�b���Aa2���O"�4ͬY/���577��Z,�%�;::BE�b1��h��/���}�A0(d�T�y�#8ΩS�~����������`w��+***22f�6
�D�T��e�L��� �tx���':::��i�4)�����]�v�s��0M�zL�wǍ��bƍ��7tt!����P(������� ��x�@��=慆��}��ǄDuuMhh�+�X�_�|���5k֋%%%MM���KS�$/]���p���{~�Q����x�"�PEE%^
�*++KNNz啅���$ɷ�:��KrGB� --�a��.�t:��Գq�����f.Z�
�0ׯ����l:����;:,���k ����{M�5D�@�j��iI�q9���H��c��%w�"���f�����F*����+0�����?���r�k[��@��^^^�� -��Egg��Y(�; ��f��{� W�Z  - h	 @K  ��  � �%  - 08P����aj��N�ˮ�	�`	H�R"��$h�qa4[[�qp2��xb(��IWҟ5Ԝ�:�Urhi�t:Z-��Ք媠a/��w��C�$�Y񯷞�?�x�4�^��}�E�$f����YtȰ���]<[#�C"J��T#��0�0��N��,h�	��y@�~i&�΁�Z(� ���BQ<��Ӄ�a-���  @K��8q�
�	���]B��g�S>�&�B���k��4�`w6B�������n��\�C�Yl���v�B�~i�^r!ю�����e����h���k2�z[���%6�5~ÓpH	�0b�8,��
]ln뤏eg�D���D"�ҥK'O�,��ZZZ*++?��S�պu�����]�v��������ϝ;�ۖcPPPrr�1c�bqNNNkkk�����eddh4��q��ŝ;w�ӆz�嗧M���x���={����-[$�瞂���Ϫ��c72<	�/��0���K]��n��{���>����oǎMMMZ�v���"��j��ڵK��?��8mڴI�&���$$$��a�A(=z�������˗��g�����������㏵�����~�5w��6@-&��j���!�+�l��H�#����o9b�1:Bl�-и�ϱ�H$JNN^�r��ӧB�/_.)��Z�d2aOpLppp|||KK˷�~�yu�F�����r�ᇛ7o����MMMB�p�ĉW�\y�XPPPPP0v�X��K��w�^�vcc�}��Z�;
�'���n-=�o��ƽ=y��S�N�����!��s�$�A�оR���#�"��DZ�p����`�A�!>ɞ�vww�4=z���ٮY�f�̙x{�����틎�NII���w;�'%%%&&FFF�ݻw�xNNNnn�����y�����7;vl{{��߿'*�*333%%[��L�����)�K��)�n�6�QȄ�ҪLH���x�?�"8N��_������_�jUff�N�;s�̱c�z����k�n߾}����E�������֭+((���G�����斔��he��������3g�4OCѿ��YYYr�\ ��/�3|5�0*�*55uĈ
�b�������|���'N��*���K4�D14��tRX�c��	�Q��W�8�s�����<xP.�oܸ������[�Fs��A��СCx���O�Ѹ�B���ø-i�=��;z��ʕ+���oll,,,<x���\�bAb�8���vǎs��]�r��ٳ��۷i�&�����y󊊊��~<#�x��3 Rσ?'�y�7UUU8Ʀ���޽{�.]�e��Q��b�� �r�!�����;ommuw�8������T\\�9ǎ�4i������G_}����zw��0����?�1,,���1jԨ�k�B�~��D8ZR�XB���(I�'�[p14ao鿪]�z����^�'�=L���e���?�N���!�@�R��Χ�����EQTIII?�2mq :233+**jjj�~?�}<��
C��f��Æ��_��j�t}p؀��t7�|��(EQ�V�r���������t�i�N������ʲ����;w�\vv6�R���m4{��ILL����>��H��Z��-����Z�Ɲ��].##kC(����>�mzz:N�R�֯____��'��>������|�D��ڙ8L�]���o���2Z�:y���a}�����3�{��r�����,Y�p8h�&I���𫯾�q�M�6��啕��4}����tnn�m���˝N��n����xc/   55u�ƍC{�)))[�n���;/_��ܹs��������X�b��͝����֭[o��fSSS�d����֭[m6�@ ���\�z5���e�'W�l6�=O�����w�h�?�ð���?��>����j5�0w���#�Ɣ F�i6�{�4��ihh��aWk��i�}nl�Yyyy�������}H&�)
���]///�Db4q<�fۛ'ʦLI��>X�o�KrFz�fs���?d��M7���ns��������0[H��[𴍑.^�x�'�����inn��詟l�a2^B�������~	ؖ��3kX�s�����qLL?�l��h�tO�ݒ��N�T�l,~�D�[��W���96=�@Kn�X,�������^��b�X,Bz��`���ү� 0^  � ����B]4GE�<@s(��A,���# �H�&E�<`��A�3|�Zz���椅cUL�9�0n���	j���R"D�e��c�fk��!NB�I3f��Ն�?XjNJ��AŌ-K����fw8i�e6\����*�BJ�ԉipPBr����E�P  Z � ��   - h	 @K  Z  � O��@a�攥u    IEND�B`�