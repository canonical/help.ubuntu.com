<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Var kan du lagra din säkerhetskopia</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#backup" title="Säkerhetskopiering">Säkerhetskopiering</a> » <a class="trail" href="backup-why.html" title="Säkerhetskopiera dina viktiga filer">Säkerhetskopior</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Var kan du lagra din säkerhetskopia</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du bör spara säkerhetskopiera av dina filer någonstans separat från din dator - till exempel på en extern hårddisk. På så sätt kan säkerhetskopia fortfarande finnas intakt om datorn går sönder. För maximal säkerhet bör du inte ha säkerhetskopia i samma byggnad som din dator. Om en brand eller inbrott inträffar så kan båda kopiorna av data gå förlorade om de lagras på samma plats.</p>
<p class="p">Det är också viktigt att välja ett lämpligt <span class="em">medium för säkerhetskopiering</span>. Du måste lagra dina säkerhetskopior på en enhet som har tillräckligt med lagringsutrymme för alla säkerhetskopierade filer.</p>
<div class="list"><div class="inner">
<div class="title title-list"><h2><span class="title">Alternativ för lokal- och fjärrlagring</span></h2></div>
<div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">USB-minne (medelkapacitet)</p></li>
<li class="list"><p class="p">Brännbar CD eller DVD (låg/medelkapacitet)</p></li>
<li class="list"><p class="p">Extern hårddisk (i regel hög kapacitet)</p></li>
<li class="list"><p class="p">Intern hårddisk (hög kapacitet)</p></li>
<li class="list"><p class="p">Nätverksansluten hårddisk (hög kapacitet)</p></li>
<li class="list"><p class="p">Fil-/säkerhetskopieringsserver (hög kapacitet)</p></li>
<li class="list"><p class="p">Säkerhetskopieringstjänst på nätet (till exempel <span class="link"><a href="http://aws.amazon.com/s3/" title="http://aws.amazon.com/s3/">Amazon S3</a></span>; kapacitet varierar efter pris)</p></li>
</ul></div>
</div></div>
<p class="p">Vissa av de här alternativen har tillräcklig kapacitet för att möjliggöra en säkerhetskopiering av alla filer på ditt system, vilket också kallas en <span class="em">fullständig systemkopiering</span>.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="backup-why.html" title="Säkerhetskopiera dina viktiga filer">Säkerhetskopiera dina viktiga filer</a><span class="desc"> — Varför, vad, var, och hur man säkerhetskopierar.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
