<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Referenser</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = "index.html.en";
        } else {
                window.location = href.replace(/\.html.*/, ".html.en");
        }
         return false;
      }
      function browserPreferredLanguage() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = href;
        } else {
                window.location = href.replace(/\.html.*/, ".html");
        }
        return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../18.04" class="trail">Ubuntu 18.04</a> » <a class="trail" href="index.html.sv" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="version-control-system.html.sv" title="Versionshanteringssystem">Versionshanteringssystem</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="subversion.html.sv" title="Subversion">Föregående</a><a class="nextlinks-next" href="samba.html.sv" title="Samba">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Referenser</h1></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
        <p class="para">
        <a href="http://bazaar.canonical.com/en/" class="ulink" title="http://bazaar.canonical.com/en/">Webbsidan för Bazaar</a>
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        <a href="https://launchpad.net/" class="ulink" title="https://launchpad.net/">Launchpad</a>
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        <a href="http://git-scm.com" class="ulink" title="http://git-scm.com">Git homepage</a>
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        <a href="https://github.com/sitaramc/gitolite" class="ulink" title="https://github.com/sitaramc/gitolite">Gitolite</a>
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        <a href="http://subversion.apache.org/" class="ulink" title="http://subversion.apache.org/">Subversions webbplats</a>
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        <a href="http://svnbook.red-bean.com/" class="ulink" title="http://svnbook.red-bean.com/">Subversion-bok</a>
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        <a href="https://help.ubuntu.com/community/EasyBazaar" class="ulink" title="https://help.ubuntu.com/community/EasyBazaar">Easy Bazaar Ubuntu Wiki page</a>
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        <a href="https://help.ubuntu.com/community/Subversion" class="ulink" title="https://help.ubuntu.com/community/Subversion">Ubuntu Wiki Subversion page</a>
        </p>
      </li>
</ul></div></div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="subversion.html.sv" title="Subversion">Föregående</a><a class="nextlinks-next" href="samba.html.sv" title="Samba">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address
          so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>
          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p>
</div>
</div>
</body>
</html>
