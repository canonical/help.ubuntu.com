<?xml version="1.0" encoding="utf-8" standalone="no"?>
<svg xmlns:osb="http://www.openswatchbook.org/uri/2009/osb" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:cc="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" xmlns:svg="http://www.w3.org/2000/svg" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" xmlns:sodipodi="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:inkscape="http://www.inkscape.org/namespaces/inkscape" height="500" id="svg10075" version="1.1" width="840" sodipodi:docname="gs-goa2.svg" inkscape:version="0.92.2 5c3e80d, 2017-08-06">
  <defs id="defs10077">
    <linearGradient id="RHEL7" osb:paint="gradient">
      <stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </linearGradient>
    <linearGradient id="GNOME" osb:paint="gradient">
      <stop id="stop11074" offset="0" style="stop-color:#eeedec;stop-opacity:1;"/>
      <stop id="stop11076" offset="1" style="stop-color:#eeedec;stop-opacity:1"/>
    </linearGradient>
    <linearGradient id="BLANK" osb:paint="gradient">
      <stop id="stop7012" offset="0" style="stop-color:#eeedec;stop-opacity:0;"/>
      <stop id="stop7014" offset="1" style="stop-color:#eeedec;stop-opacity:0"/>
    </linearGradient>
    <linearGradient gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" gradientUnits="userSpaceOnUse" id="linearGradient7064" x1="-18.33782" x2="713.42853" y1="490.54935" y2="490.54935" inkscape:collect="always" xlink:href="#GNOME"/>
    <filter color-interpolation-filters="sRGB" height="1.1308649" id="filter5601" width="1.2058235" x="-0.10291173" y="-0.065432459" inkscape:collect="always">
      <feGaussianBlur id="feGaussianBlur5603" stdDeviation="0.610872" inkscape:collect="always"/>
    </filter>
    <linearGradient gradientUnits="userSpaceOnUse" id="linearGradient5885" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" inkscape:collect="always" xlink:href="#linearGradient5716"/>
    <linearGradient id="linearGradient5716">
      <stop id="stop5718" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <stop id="stop5720" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </linearGradient>
    <linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17441" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" inkscape:collect="always" xlink:href="#linearGradient5716"/>
    <linearGradient id="linearGradient17443">
      <stop id="stop17445" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <stop id="stop17447" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </linearGradient>
    <linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17453" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" inkscape:collect="always" xlink:href="#linearGradient5716"/>
    <linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17455" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" inkscape:collect="always" xlink:href="#linearGradient5716"/>
  </defs>
  <sodipodi:namedview bordercolor="#666666" borderlayer="true" borderopacity="1.0" fit-margin-bottom="0" fit-margin-left="0" fit-margin-right="0" fit-margin-top="0" height="0px" id="base" pagecolor="#eeeeec" showgrid="false" width="0px" inkscape:current-layer="g4890" inkscape:cx="244.2324" inkscape:cy="43.939731" inkscape:document-units="px" inkscape:pageopacity="1" inkscape:pageshadow="2" inkscape:showpageshadow="false" inkscape:window-height="1403" inkscape:window-maximized="1" inkscape:window-width="2560" inkscape:window-x="3440" inkscape:window-y="0" inkscape:zoom="1" inkscape:document-rotation="0">
    <inkscape:grid empspacing="5" enabled="true" id="grid17504" snapvisiblegridlinesonly="true" type="xygrid" visible="true"/>
  </sodipodi:namedview>
  <metadata id="metadata10080">
    <rdf:RDF>
      <cc:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </cc:Work>
    </rdf:RDF>
  </metadata>
  <g id="layer1" transform="translate(0,-992.3622)" sodipodi:insensitive="true" inkscape:groupmode="layer" inkscape:label="bg">
    <rect height="656" id="background" style="fill:url(#BLANK);" width="866" x="-16" y="855.36218" inkscape:label="background"/>
  </g>
  <g id="layer2" transform="translate(0,-540)" inkscape:groupmode="layer" inkscape:label="fg">
    <g id="g11020" transform="translate(-35,-139.36217)">
      <path d="m 137,278 a 17,17 0 0 1 -17,17 17,17 0 0 1 -17,-17 17,17 0 0 1 17,-17 17,17 0 0 1 17,17 z" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(2,453.36217)" sodipodi:cx="120" sodipodi:cy="278" sodipodi:rx="17" sodipodi:ry="17" sodipodi:type="arc"/>
      <text id="text11016" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" xml:space="preserve"><tspan id="tspan11018" x="122.29289" y="736.36218" sodipodi:role="line" style="font-size:14px;line-height:1.25">3</tspan></text>
    </g>
    <g id="g4890" style="display:inline" transform="matrix(2.6833333,0,0,2.6833333,-1275.5101,-1072.8539)">
      <path d="m 528.04724,634.48596 h 209.13044 c 2.216,0 4,1.7996 4,4.03497 v 122.79112 h -4 -209.13044 -4 V 638.52093 c 0,-2.23537 1.784,-4.03497 4,-4.03497 z" id="path5430" style="fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-opacity:1" sodipodi:nodetypes="sssccccss" inkscape:connector-curvature="0"/>
      <path d="m 524.59833,653.09463 c 212.46132,0 216.29809,0 216.29809,0" id="path5361" style="fill:none;stroke:#000000;stroke-width:1.01455009;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" inkscape:connector-curvature="0"/>
      <g id="g5363" style="fill:#0c0000;fill-opacity:1" transform="matrix(0.47058484,0,0,0.47058484,728.13789,640.56125)">
        <g id="g5365" style="display:inline;fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5367" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5369" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5371" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)">
          <g id="g5373" style="display:inline;fill:#0c0000;fill-opacity:1" transform="translate(19,-242)">
            <path d="m 45,764 h 1 c 0.01037,-1.2e-4 0.02079,-4.6e-4 0.03125,0 0.254951,0.0112 0.50987,0.12858 0.6875,0.3125 L 49,766.59375 51.3125,764.3125 C 51.578125,764.082 51.759172,764.007 52,764 h 1 v 1 c 0,0.28647 -0.03434,0.55065 -0.25,0.75 l -2.28125,2.28125 2.25,2.25 C 52.906938,770.46942 52.999992,770.7347 53,771 v 1 h -1 c -0.265301,-10e-6 -0.530586,-0.0931 -0.71875,-0.28125 L 49,769.4375 46.71875,771.71875 C 46.530586,771.90694 46.26529,772 46,772 h -1 v -1 c -3e-6,-0.26529 0.09306,-0.53058 0.28125,-0.71875 l 2.28125,-2.25 L 45.28125,765.75 C 45.070508,765.55537 44.97809,765.28075 45,765 Z" id="path5375" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.78124988;marker:none;enable-background:new" inkscape:connector-curvature="0"/>
          </g>
        </g>
        <g id="g5377" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5379" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5381" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
      </g>
      <text id="text12012" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none" x="634.84845" y="645.41119" xml:space="preserve"><tspan id="tspan12014" x="634.84845" y="645.41119" sodipodi:role="line" style="font-size:5.21739101px;line-height:1.25">Nätkonton</tspan></text>
      <rect style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:0.37267083;stroke-opacity:1" id="rect884" width="180.65475" height="63.068722" x="546.07709" y="698.2431"/>
      <g id="default-pointer-c" style="display:inline" transform="matrix(1.0281734,0,0,1.0281734,656.14965,720.60298)" inkscape:label="#g5607">
        <path d="M 27.135224,2.8483222 V 19.288556 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path5567" style="color:#000000;display:block;overflow:visible;visibility:visible;opacity:0.6;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;filter:url(#filter5601);enable-background:accumulate" sodipodi:nodetypes="cccccccc" inkscape:connector-curvature="0"/>
        <path d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path5565" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17453);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" sodipodi:nodetypes="cccccccc" inkscape:connector-curvature="0"/>
        <path d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path6242" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17455);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" sodipodi:nodetypes="cccccccc" inkscape:connector-curvature="0"/>
      </g>
      <g id="g4705" style="display:inline" transform="matrix(0.37267081,0,0,0.37267081,492.83185,447.51482)" inkscape:label="go-previous">
        <rect height="16" id="rect10837-5-8-1" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none;enable-background:new" transform="scale(-1,1)" width="16" x="-116" y="518"/>
        <path d="m 112.01352,520 h -1 c -0.0104,-1.2e-4 -0.0208,-4.6e-4 -0.0313,0 -0.25495,0.0112 -0.50987,0.12858 -0.6875,0.3125 l -6.29767,5.71875 6.29772,5.71875 c 0.18816,0.18819 0.45346,0.28125 0.71875,0.28125 h 1 v -1 c 0,-0.26529 -0.0931,-0.53058 -0.28125,-0.71875 l -4.82897,-4.28125 4.82897,-4.28125 c 0.21074,-0.19463 0.30316,-0.46925 0.28125,-0.75 z" id="path10839-9-9-5" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.78124988;marker:none;enable-background:new" sodipodi:nodetypes="ccsccccccccccc" inkscape:connector-curvature="0"/>
      </g>
      <rect height="11.925466" id="rect15386" rx="1.4906832" ry="1.4906832" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.3726708;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" width="11.925466" x="527.34424" y="637.76007"/>
      <rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:7.45341635;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect977" width="2.6351805" height="45.325108" x="734.86548" y="657.14594" rx="1.3175902" ry="1.3175902"/>
      <rect y="705.88513" x="555.11969" height="14.863034" width="15.262931" id="rect979" style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:0.37267083;stroke-opacity:1"/>
      <rect style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:0.37267083;stroke-opacity:1" id="rect981" width="15.262931" height="14.863034" x="555.11969" y="728.24542"/>
      <rect y="750.60571" x="555.11969" height="10.70611" width="15.262931" id="rect983" style="color:#000000;overflow:visible;opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:0.37267083;stroke-opacity:1"/>
      <rect style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:7.45341635;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect985" width="66.406548" height="7.3785057" x="576.00928" y="709.38965"/>
      <rect y="731.26166" x="576.00928" height="7.3785057" width="47.433247" id="rect987" style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:7.45341635;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal"/>
      <rect style="opacity:1;vector-effect:none;fill:#d3d7cf;fill-opacity:1;stroke:none;stroke-width:7.45341635;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect989" width="75.893196" height="5.392509" x="576.00928" y="753.66071"/>
      <flowRoot xml:space="preserve" id="flowRoot1005" style="fill:black;fill-opacity:1;stroke:none;font-family:sans-serif;font-style:normal;font-weight:normal;font-size:40px;line-height:1.25;letter-spacing:0px;word-spacing:0px"><flowRegion id="flowRegion1007"><rect id="rect1009" width="488" height="122" x="186" y="199"/></flowRegion><flowPara id="flowPara1011"/></flowRoot>      <text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.46583891px;line-height:1.25;font-family:sans-serif;-inkscape-font-specification:'sans-serif, Normal';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" x="546.89825" y="693.11334" id="text1074"><tspan sodipodi:role="line" id="tspan1072" x="546.89825" y="693.11334" style="stroke-width:0.3726708">Add an account</tspan></text>
      <g id="g3922" style="display:inline;stroke-width:0.80000001" transform="matrix(0.93167703,0,0,0.93167703,417.23142,562.40689)" inkscape:label="account-facebook">
        <rect height="16" id="rect2941" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.80000001;marker:none" transform="rotate(-90)" width="16" x="-194" y="20" inkscape:label="audio-volume-high"/>
        <path d="M 22.116732,178 C 20.946094,178 20,178.94979 20,180.125 v 11.75 c 0,1.17521 0.946094,2.125 2.116732,2.125 h 6.910506 v -6 h -0.99611 v -2 h 0.99611 v -1.0625 c 0,-1.84445 1.374066,-2.88912 3.175096,-2.9375 h 1.77432 v 2 H 32.88716 c -0.625856,0 -0.902724,0.22291 -0.902724,0.90625 V 186 h 1.712062 l -0.217898,2 h -1.494164 v 6 h 1.898832 C 35.053906,194 36,193.05021 36,191.875 v -11.75 C 36,178.94979 35.053906,178 33.883268,178 Z" id="rect14063" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.40000001;marker:none;enable-background:new" sodipodi:nodetypes="sssscccccscccsscccccsssss" inkscape:connector-curvature="0"/>
      </g>
      <path d="m 440.17988,706.63884 -1.65949,-0.006 c -1.16975,0.60941 -1.34475,2.13001 -0.96077,3.52277 0.50753,1.84074 1.52186,3.13191 2.88229,2.70761 1.89768,-0.59201 1.95321,-2.14178 1.36835,-3.95949 -0.30932,-0.9614 -0.88305,-1.73598 -1.63038,-2.26361 z m 4.62912,2.87499 c 0,0.81962 -0.33349,1.51919 -0.69873,2.06709 v 0.0293 l -0.0874,0.0582 c 0,0 -0.23734,0.27876 -0.52405,0.55318 -0.2863,0.27447 -0.72785,0.64051 -0.72785,0.64051 -0.35929,0.27003 -0.55315,0.627 -0.55315,1.01897 0,0.39332 0.24992,0.74883 0.61139,1.01899 0,0 0.73301,0.44913 1.13544,0.78609 0.40226,0.33716 0.87343,0.78607 0.87343,0.78607 0.54483,0.51229 0.90252,1.32866 0.90252,2.24177 0,0.78641 -0.24936,1.49952 -0.66962,2.00886 l -0.64051,0.8152 h 3.9886 c 1.09064,0 1.97976,-0.88488 1.97976,-1.97976 v -10.94684 c 0,-1.09487 -0.88912,-1.97974 -1.97976,-1.97974 -0.53462,-0.005 -1.69697,10e-4 -1.69697,10e-4 l -0.0143,0.91826 -2.39058,0.26813 c 0.3498,0.60748 0.4829,1.21381 0.49188,1.69431 z m -9.31647,2.2709 v 5.2405 c 1.61776,-1.08314 4.51267,-1.10633 4.51267,-1.10633 0,0 0.0125,-0.0175 0,-0.0293 -1.16064,-0.89223 -0.66962,-1.92158 -0.66962,-1.92158 -1.79456,0.15289 -2.61487,-0.51693 -3.84305,-2.18353 z m 4.71648,5.15317 c -1.61229,0.0906 -3.68685,0.75809 -3.72659,2.35822 0,0.95714 0.6231,1.82472 1.51391,2.21266 0,0 0.032,0.0205 0.0582,0.0293 h 0.0293 4.22152 c 0,0 0.008,-0.0417 0.0293,-0.0582 2.28366,-2.0211 0.55915,-3.19293 -1.39748,-4.51265 -0.0355,-0.0236 -0.0874,-0.0293 -0.0874,-0.0293 -0.20403,-0.008 -0.41019,-0.0128 -0.6405,0 z" id="path14750" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.1863354;marker:none;enable-background:new" sodipodi:nodetypes="ccccscscccccscccsccssscccccsccccsccccccccsccc" inkscape:connector-curvature="0"/>
    </g>
    <text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:21.33333397px;line-height:1.25;font-family:sans-serif;-inkscape-font-specification:'sans-serif, Normal';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1" x="420" y="735" id="text1050"><tspan sodipodi:role="line" id="tspan1048" x="420" y="735">Connect to your data in the cloud</tspan></text>
  </g>
</svg>
