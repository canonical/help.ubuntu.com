<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Filer, mappar och sökning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 25.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Filer, mappar och sökning</span></h1></div>
<div class="region">
<div class="contents pagewide"></div>
<section id="common-file-tasks"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Vanliga åtgärder</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="files-browse.html.sv" title="Bläddra bland filer och mappar"><span class="title">Bläddra bland filer och mappar</span><span class="linkdiv-dash"> — </span><span class="desc">Hantera och organisera filer med filhanteraren.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-rename.html.sv" title="Byt namn på en fil eller mapp"><span class="title">Byt namn på en fil eller mapp</span><span class="linkdiv-dash"> — </span><span class="desc">Byt namn på fil eller mapp.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-rename-multiple.html.sv" title="Byt namn på flera filer"><span class="title">Byt namn på flera filer</span><span class="linkdiv-dash"> — </span><span class="desc">Byt namn på mer än en fil samtidigt.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-rename-music-metadata.html.sv" title="Byt namn på musikfiler med hjälp av metadata"><span class="title">Byt namn på musikfiler med hjälp av metadata</span><span class="linkdiv-dash"> — </span><span class="desc">Byt namn på musikfiler med hjälp av metadata de innehåller.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-preview.html.sv" title="Förhandsgranska filer och mappar"><span class="title">Förhandsgranska filer och mappar</span><span class="linkdiv-dash"> — </span><span class="desc">Visa och dölj snabbt förhandsgranskningar av dokument, bilder, videor och mera.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="files-copy.html.sv" title="Kopiera eller flytta filer och mappar"><span class="title">Kopiera eller flytta filer och mappar</span><span class="linkdiv-dash"> — </span><span class="desc">Kopiera eller flytta objekt till en ny mapp.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-sort.html.sv" title="Sortera filer och mappar"><span class="title">Sortera filer och mappar</span><span class="linkdiv-dash"> — </span><span class="desc">Sortera filer efter namn, storlek, typ, eller när de ändrades.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-search.html.sv" title="Sök efter filer"><span class="title">Sök efter filer</span><span class="linkdiv-dash"> — </span><span class="desc">Hitta filer baserat på filnamn och typ.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-delete.html.sv" title="Ta bort filer och mappar"><span class="title">Ta bort filer och mappar</span><span class="linkdiv-dash"> — </span><span class="desc">Ta bort filer eller mappar som du inte längre behöver.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="more-file-tasks"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Fler filrelaterade uppgifter</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="nautilus-connect.html.sv" title="Bläddra genom filer på en server eller nätverksutdelning"><span class="title">Bläddra genom filer på en server eller nätverksutdelning</span><span class="linkdiv-dash"> — </span><span class="desc">Titta på och redigera filer på en annan dator över FTP, SSH, Windows-utdelningar eller WebDAV.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-share.html.sv" title="Dela filer visa e-post"><span class="title">Dela filer visa e-post</span><span class="linkdiv-dash"> — </span><span class="desc">Överför enkelt filer till dina e-postkontakter från filhanteraren.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="nautilus-file-properties-basic.html.sv" title="Filegenskaper"><span class="title">Filegenskaper</span><span class="linkdiv-dash"> — </span><span class="desc">Visa grundläggande filinformation, ställa in rättigheter och välja standardprogram.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-lost.html.sv" title="Hitta en borttappad fil"><span class="title">Hitta en borttappad fil</span><span class="linkdiv-dash"> — </span><span class="desc">Följ dessa tips om du inte kan hitta en fil du har skapat eller hämtat.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="nautilus-prefs.html.sv" title="Inställningar för filhanterare"><span class="title">Inställningar för filhanterare</span><span class="linkdiv-dash"> — </span><span class="desc">Visa och ställ in inställningar för filhanteraren.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="files-disc-write.html.sv" title="Skriv filer till en cd- eller dvd-skiva"><span class="title">Skriv filer till en cd- eller dvd-skiva</span><span class="linkdiv-dash"> — </span><span class="desc">Spara undan filer och dokument på en blank cd eller dvd med hjälp av en cd/dvd-brännare.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="privacy-history-recent-off.html.sv" title="Stäng av eller begränsa filhistorik"><span class="title">Stäng av eller begränsa filhistorik</span><span class="linkdiv-dash"> — </span><span class="desc">Stoppa eller begränsa din dator från att spåra dina nyligen använda filer.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="privacy-purge.html.sv" title="Töm papperskorgen &amp; ta bort tillfälliga filer"><span class="title">Töm papperskorgen &amp; ta bort tillfälliga filer</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in hur ofta din papperskorg och tillfälliga filer kommer att rensas bort från din dator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-recover.html.sv" title="Återskapa en fil från Papperskorgen"><span class="title">Återskapa en fil från Papperskorgen</span><span class="linkdiv-dash"> — </span><span class="desc">Borttagna filer skickas normalt till Papperskorgen, men kan återställas.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-open.html.sv" title="Öppna filer med andra program"><span class="title">Öppna filer med andra program</span><span class="linkdiv-dash"> — </span><span class="desc">Öppna filer med ett program som inte är standardprogrammet för den typen av fil. Du kan även ändra standardprogrammet.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="removable"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Flyttbara enheter och externa diskar</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs"><div class="linkdiv "><a class="linkdiv" href="files-removedrive.html.sv" title="Säker borttagning av extern enhet"><span class="title">Säker borttagning av extern enhet</span><span class="linkdiv-dash"> — </span><span class="desc">Mata ut eller avmontera en USB-enhet, cd, dvd eller annan enhet.</span></a></div></div>
<div class="links-divs"><div class="linkdiv "><a class="linkdiv" href="files-autorun.html.sv" title="Öppna program för enheter eller diskar"><span class="title">Öppna program för enheter eller diskar</span><span class="linkdiv-dash"> — </span><span class="desc">Kör automatiskt program för cd och dvd, kameror, musikspelare, och andra enheter och media.</span></a></div></div>
</div></div></div></div></div></div>
</div></section><section id="backup"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Säkerhetskopiering</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="backup-frequency.html.sv" title="Frekvens för säkerhetskopiering"><span class="title">Frekvens för säkerhetskopiering</span><span class="linkdiv-dash"> — </span><span class="desc">Lär dig hur ofta du bör säkerhetskopiera dina viktiga filer för att se till att de är säkra.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="backup-check.html.sv" title="Kontrollera din säkerhetskopia"><span class="title">Kontrollera din säkerhetskopia</span><span class="linkdiv-dash"> — </span><span class="desc">Verifiera att din säkerhetskopiering lyckades.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="backup-why.html.sv" title="Säkerhetskopiera dina viktiga filer"><span class="title">Säkerhetskopiera dina viktiga filer</span><span class="linkdiv-dash"> — </span><span class="desc">Varför, vad, var och hur man säkerhetskopierar.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="backup-thinkabout.html.sv" title="Var kan jag hitta filerna jag vill säkerhetskopiera?"><span class="title">Var kan jag hitta filerna jag vill säkerhetskopiera?</span><span class="linkdiv-dash"> — </span><span class="desc">En lista över mappar där du kan hitta dokument, filer och inställningar som du kanske vill säkerhetskopiera.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="backup-restore.html.sv" title="Återställ en säkerhetskopia"><span class="title">Återställ en säkerhetskopia</span><span class="linkdiv-dash"> — </span><span class="desc">Återskapa dina filer från en säkerhetskopia.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="faq"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Tips och frågor</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="nautilus-file-properties-permissions.html.sv" title="Ange filrättigheter"><span class="title">Ange filrättigheter</span><span class="linkdiv-dash"> — </span><span class="desc">Styr vem som kan titta på och redigera dina filer och mappar.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-hidden.html.sv" title="Dölj en fil"><span class="title">Dölj en fil</span><span class="linkdiv-dash"> — </span><span class="desc">Gör en fil osynlig så att du inte kan se den i filhanteraren.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-templates.html.sv" title="Mallar för vanliga dokumenttyper"><span class="title">Mallar för vanliga dokumenttyper</span><span class="linkdiv-dash"> — </span><span class="desc">Skapa snabbt dokument från anpassade filmallar.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="files-select.html.sv" title="Markera filer efter mönster"><span class="title">Markera filer efter mönster</span><span class="linkdiv-dash"> — </span><span class="desc">Tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>S</kbd></span></span> för att markera flera filer som har liknande namn.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="nautilus-bookmarks-edit.html.sv" title="Redigera bokmärken för mappar"><span class="title">Redigera bokmärken för mappar</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till, ta bort och byt namn på bokmärken i filhanteraren.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-tilde.html.sv" title="Vad är en fil med en ~ i slutet på namnet?"><span class="title">Vad är en fil med en <span class="file">~</span> i slutet på namnet?</span><span class="linkdiv-dash"> — </span><span class="desc">Detta är säkerhetskopior. De är dolda som standard.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
