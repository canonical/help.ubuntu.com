<?xml version="1.0" encoding="utf-8" standalone="no"?>
<svg xmlns:osb="http://www.openswatchbook.org/uri/2009/osb" xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:cc="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" xmlns:svg="http://www.w3.org/2000/svg" xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" xmlns:sodipodi="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:inkscape="http://www.inkscape.org/namespaces/inkscape" height="1000" id="svg10075" version="1.1" width="840" sodipodi:docname="gs-goa4.svg" inkscape:version="0.92.2 5c3e80d, 2017-08-06">
  <defs id="defs10077">
    <linearGradient id="RHEL7" osb:paint="gradient">
      <stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </linearGradient>
    <linearGradient id="GNOME" osb:paint="gradient">
      <stop id="stop11074" offset="0" style="stop-color:#eeedec;stop-opacity:1;"/>
      <stop id="stop11076" offset="1" style="stop-color:#eeedec;stop-opacity:1"/>
    </linearGradient>
    <linearGradient id="BLANK" osb:paint="gradient">
      <stop id="stop7012" offset="0" style="stop-color:#eeedec;stop-opacity:0;"/>
      <stop id="stop7014" offset="1" style="stop-color:#eeedec;stop-opacity:0"/>
    </linearGradient>
    <linearGradient gradientTransform="matrix(1.1834379,0,0,1.4157524,5.7016703,-219.13426)" gradientUnits="userSpaceOnUse" id="linearGradient7064" x1="-18.33782" x2="713.42853" y1="490.54935" y2="490.54935" inkscape:collect="always" xlink:href="#GNOME"/>
    <linearGradient gradientUnits="userSpaceOnUse" id="linearGradient5885" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" inkscape:collect="always" xlink:href="#linearGradient5716"/>
    <linearGradient id="linearGradient5716">
      <stop id="stop5718" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <stop id="stop5720" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </linearGradient>
    <linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17441" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" inkscape:collect="always" xlink:href="#linearGradient5716"/>
    <linearGradient id="linearGradient17443">
      <stop id="stop17445" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <stop id="stop17447" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </linearGradient>
    <clipPath clipPathUnits="userSpaceOnUse" id="clipPath24278">
      <path d="m 0,0 0,2482 2306,0 L 2306,0 0,0 z" id="path24280" inkscape:connector-curvature="0"/>
    </clipPath>
  </defs>
  <sodipodi:namedview bordercolor="#666666" borderlayer="true" borderopacity="1.0" fit-margin-bottom="0" fit-margin-left="0" fit-margin-right="0" fit-margin-top="0" height="0px" id="base" pagecolor="#eeeeec" showgrid="false" width="0px" inkscape:current-layer="layer2" inkscape:cx="192.59471" inkscape:cy="671.89139" inkscape:document-units="px" inkscape:pageopacity="1" inkscape:pageshadow="2" inkscape:showpageshadow="false" inkscape:snap-bbox="true" inkscape:snap-nodes="false" inkscape:window-height="1403" inkscape:window-maximized="1" inkscape:window-width="2560" inkscape:window-x="3440" inkscape:window-y="0" inkscape:zoom="1">
    <inkscape:grid empspacing="5" enabled="true" id="grid17504" snapvisiblegridlinesonly="true" type="xygrid" visible="true"/>
  </sodipodi:namedview>
  <metadata id="metadata10080">
    <rdf:RDF>
      <cc:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </cc:Work>
    </rdf:RDF>
  </metadata>
  <g id="layer1" transform="translate(0,-492.3622)" sodipodi:insensitive="true" inkscape:groupmode="layer" inkscape:label="bg">
    <rect height="1036" id="background" style="fill:url(#BLANK);" width="866" x="-16" y="475.36218" inkscape:label="background"/>
    <path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:5.36666679;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" d="m 176.5,555.3622 h 487 c 9.972,0 18,8.028 18,18 v 352 h -523 v -352 c 0,-9.972 8.028,-18 18,-18 z" id="rect24979-0" inkscape:connector-curvature="0" sodipodi:nodetypes="sssccss"/>
    <text id="text24981-9" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="426.95731" y="581.19922" xml:space="preserve"><tspan id="tspan24983-4" x="426.95731" y="581.19922" sodipodi:role="line" style="font-size:14px;line-height:1.25">Google-konto</tspan></text>
    <g id="g5363-3" style="display:inline;fill:#0c0000;fill-opacity:1" transform="matrix(1.262736,0,0,1.262736,644.9001,569.2605)">
      <g id="g5365-3" style="display:inline;fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
      <g id="g5367-2" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
      <g id="g5369-7" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
      <g id="g5371-9" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)">
        <g id="g5373-7" style="display:inline;fill:#0c0000;fill-opacity:1" transform="translate(19,-242)">
          <path d="m 45,764 h 1 c 0.01037,-1.2e-4 0.02079,-4.6e-4 0.03125,0 0.254951,0.0112 0.50987,0.12858 0.6875,0.3125 L 49,766.59375 51.3125,764.3125 C 51.578125,764.082 51.759172,764.007 52,764 h 1 v 1 c 0,0.28647 -0.03434,0.55065 -0.25,0.75 l -2.28125,2.28125 2.25,2.25 C 52.906938,770.46942 52.999992,770.7347 53,771 v 1 h -1 c -0.265301,-10e-6 -0.530586,-0.0931 -0.71875,-0.28125 L 49,769.4375 46.71875,771.71875 C 46.530586,771.90694 46.26529,772 46,772 h -1 v -1 c -3e-6,-0.26529 0.09306,-0.53058 0.28125,-0.71875 l 2.28125,-2.25 L 45.28125,765.75 C 45.070508,765.55537 44.97809,765.28075 45,765 Z" id="path5375-1" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.78124988;marker:none;enable-background:new" inkscape:connector-curvature="0"/>
        </g>
      </g>
      <g id="g5377-8" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
      <g id="g5379-9" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
      <g id="g5381-5" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
    </g>
  </g>
  <g id="layer2" transform="translate(0,-40)" inkscape:groupmode="layer" inkscape:label="fg">
    <g id="g11020" transform="translate(-35,-619.36217)">
      <path d="m 137,278 a 17,17 0 0 1 -17,17 17,17 0 0 1 -17,-17 17,17 0 0 1 17,-17 17,17 0 0 1 17,17 z" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(2,453.36217)" sodipodi:cx="120" sodipodi:cy="278" sodipodi:rx="17" sodipodi:ry="17" sodipodi:type="arc"/>
      <text id="text11016" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" xml:space="preserve"><tspan id="tspan11018" x="122.29289" y="736.36218" sodipodi:role="line" style="font-size:14px;line-height:1.25">5</tspan></text>
    </g>
    <rect y="150" x="167.50003" width="505.19278" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#eeeeec;stroke:#000000;stroke-width:1.96981525;stroke-opacity:1;marker:none;enable-background:accumulate" ry="0.36744055" rx="0.38461545" id="rect12010-4" height="313.93021"/>
    <text xml:space="preserve" y="206" x="180.5" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:sans-serif;-inkscape-font-specification:Sans;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" id="text24901"><tspan style="font-size:14px;line-height:1.25;font-family:sans-serif" sodipodi:role="line" y="206" x="180.5" id="tspan24903">Logga in</tspan></text>
    <text xml:space="preserve" y="239" x="180.5" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:sans-serif;-inkscape-font-specification:'Sans Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" id="text24905"><tspan style="font-size:13px;line-height:1.25;font-family:sans-serif" sodipodi:role="line" y="239" x="180.5" id="tspan24907">E-post</tspan></text>
    <rect y="245.5" x="182" width="480" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#babdb6;stroke-width:1;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" ry="0.36744055" rx="0.38461545" id="rect24909" height="35"/>
    <text xml:space="preserve" y="309" x="180.5" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:sans-serif;-inkscape-font-specification:'Sans Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" id="text24911"><tspan style="font-size:13px;line-height:1.25;font-family:sans-serif" sodipodi:role="line" y="309" x="180.5" id="tspan24913">Lösenord</tspan></text>
    <rect y="315.5" x="182" width="480" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#babdb6;stroke-width:1;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" ry="0.36744055" rx="0.38461545" id="rect24915" height="35"/>
    <rect y="365" x="181.5" width="106" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#729fcf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" id="rect24917" height="34"/>
    <text xml:space="preserve" y="386" x="235.5" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" id="text24919"><tspan style="font-size:12px;line-height:1.25" sodipodi:role="line" y="386" x="235.5" id="tspan24921">Logga in</tspan></text>
    <text xml:space="preserve" y="267" x="190.5" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:sans-serif;-inkscape-font-specification:Sans;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" id="text24923"><tspan style="font-size:14px;line-height:1.25;font-family:sans-serif" sodipodi:role="line" y="267" x="190.5" id="tspan24925">maria.johansson@gmail.com</tspan></text>
    <circle r="6.5" cy="332.5" cx="198" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;enable-background:accumulate" id="path24927"/>
    <circle r="6.5" cy="332.5" cx="214" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;enable-background:accumulate" id="path24929"/>
    <circle r="6.5" cy="332.5" cx="230" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;enable-background:accumulate" id="path24931"/>
    <circle r="6.5" cy="332.5" cx="246" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;enable-background:accumulate" id="path24933"/>
    <circle r="6.5" cy="332.5" cx="262" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;enable-background:accumulate" id="path24935"/>
    <g id="g24977" transform="translate(17.5,460)">
      <path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:5.36666679;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" d="m 159,105 h 487 c 9.972,0 18,8.028 18,18 v 351.99997 l -523,0 V 123 c 0,-9.972 8.028,-18 18,-18 z" id="rect24979" inkscape:connector-curvature="0" sodipodi:nodetypes="sssccss"/>
      <text id="text24981" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="409.45731" y="130.83698" xml:space="preserve"><tspan id="tspan24983" x="409.45731" y="130.83698" sodipodi:role="line" style="font-size:14px;line-height:1.25">Google-konto</tspan></text>
      <rect height="313.93021" id="rect24985" rx="0.38461545" ry="0.36744055" style="color:#000000;fill:#eeeeec;stroke:#000000;stroke-width:1.96981525;stroke-opacity:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="505.19278" x="150.00003" y="150"/>
      <rect height="16" id="rect25076" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="451" x="164" y="167"/>
      <rect height="16" id="rect25078" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="274" x="164" y="192"/>
      <rect height="16" id="rect25085" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="119" x="164" y="231"/>
      <rect height="16" id="rect25087" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="95" x="164" y="256"/>
      <rect height="16" id="rect25089" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="119" x="164" y="281"/>
      <rect height="16" id="rect25091" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="95" x="164" y="306"/>
      <rect height="311" id="rect25093" style="color:#000000;fill:#d3d7cf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="16" x="638.5" y="151"/>
      <rect height="203" id="rect25095" rx="4.1756759" ry="4.1756759" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#888a85;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="8.3513517" x="642.5" y="252"/>
      <g id="g5363" style="display:inline;fill:#0c0000;fill-opacity:1" transform="matrix(1.262736,0,0,1.262736,627.4001,118.89826)">
        <g id="g5365" style="display:inline;fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5367" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5369" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5371" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)">
          <g id="g5373" style="display:inline;fill:#0c0000;fill-opacity:1" transform="translate(19,-242)">
            <path d="m 45,764 h 1 c 0.01037,-1.2e-4 0.02079,-4.6e-4 0.03125,0 0.254951,0.0112 0.50987,0.12858 0.6875,0.3125 L 49,766.59375 51.3125,764.3125 C 51.578125,764.082 51.759172,764.007 52,764 h 1 v 1 c 0,0.28647 -0.03434,0.55065 -0.25,0.75 l -2.28125,2.28125 2.25,2.25 C 52.906938,770.46942 52.999992,770.7347 53,771 v 1 h -1 c -0.265301,-10e-6 -0.530586,-0.0931 -0.71875,-0.28125 L 49,769.4375 46.71875,771.71875 C 46.530586,771.90694 46.26529,772 46,772 h -1 v -1 c -3e-6,-0.26529 0.09306,-0.53058 0.28125,-0.71875 l 2.28125,-2.25 L 45.28125,765.75 C 45.070508,765.55537 44.97809,765.28075 45,765 Z" id="path5375" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.78124988;marker:none;enable-background:new" inkscape:connector-curvature="0"/>
          </g>
        </g>
        <g id="g5377" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5379" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
        <g id="g5381" style="fill:#0c0000;fill-opacity:1" transform="translate(-60,-518)"/>
      </g>
    </g>
    <g id="g25055" transform="translate(-35,-159.36217)">
      <path d="m 137,278 a 17,17 0 0 1 -17,17 17,17 0 0 1 -17,-17 17,17 0 0 1 17,-17 17,17 0 0 1 17,17 z" id="path25057" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(2,453.36217)" sodipodi:cx="120" sodipodi:cy="278" sodipodi:rx="17" sodipodi:ry="17" sodipodi:type="arc"/>
      <text id="text25059" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" xml:space="preserve"><tspan id="tspan25061" x="122.29289" y="736.36218" sodipodi:role="line" style="font-size:14px;line-height:1.25">6</tspan></text>
    </g>
    <rect height="34" id="rect24917-8" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#729fcf;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:5.36666679;marker:none;enable-background:accumulate" width="106" x="527" y="861" rx="8" ry="8"/>
    <text id="text24919-8" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="581" y="882" xml:space="preserve"><tspan id="tspan24921-0" x="581" y="882" sodipodi:role="line" style="font-size:12px;line-height:1.25">ALLOW</tspan></text>
    <text xml:space="preserve" y="882" x="461" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#729fcf;fill-opacity:1;stroke:none" id="text3888"><tspan style="font-size:12px;line-height:1.25;fill:#729fcf;fill-opacity:1" sodipodi:role="line" y="882" x="461" id="tspan3886">CANCEL</tspan></text>
  </g>
  <g id="layer3" style="display:none" inkscape:groupmode="layer" inkscape:label="stuff">
    <text id="text17640" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="-218.54269" y="669.83698" xml:space="preserve"><tspan id="tspan17642" x="-218.54269" y="669.83698" sodipodi:role="line" style="font-size:14px;line-height:1.25">Google</tspan></text>
    <text id="text17893" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="-218.54269" y="709.83698" xml:space="preserve"><tspan id="tspan17895" x="-218.54269" y="709.83698" sodipodi:role="line" style="font-size:14px;line-height:1.25">Facebook</tspan></text>
    <text id="text17897" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="-218.54269" y="749.83698" xml:space="preserve"><tspan id="tspan17899" x="-218.54269" y="749.83698" sodipodi:role="line" style="font-size:14px;line-height:1.25">Windows Live</tspan></text>
    <text id="text17901" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="-218.54269" y="789.83698" xml:space="preserve"><tspan id="tspan17903" x="-218.54269" y="789.83698" sodipodi:role="line" style="font-size:14px;line-height:1.25">Microsoft Exchange</tspan></text>
    <text id="text17905" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="-218.54269" y="829.83698" xml:space="preserve"><tspan id="tspan17907" x="-218.54269" y="829.83698" sodipodi:role="line" style="font-size:14px;line-height:1.25">Företagsinloggning (Kerberos)</tspan></text>
    <g id="g3922" style="display:inline" transform="matrix(2,0,0,2,-302,333)" inkscape:label="account-facebook">
      <rect height="16" id="rect2941" style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" transform="matrix(0,-1,1,0,0,0)" width="16" x="-194" y="20" inkscape:label="audio-volume-high"/>
      <path d="M 22.116732,178 C 20.946094,178 20,178.94979 20,180.125 l 0,11.75 c 0,1.17521 0.946094,2.125 2.116732,2.125 l 6.910506,0 0,-6 -0.99611,0 0,-2 0.99611,0 0,-1.0625 c 0,-1.84445 1.374066,-2.88912 3.175096,-2.9375 l 1.77432,0 0,2 -1.089494,0 c -0.625856,0 -0.902724,0.22291 -0.902724,0.90625 l 0,1.09375 1.712062,0 -0.217898,2 -1.494164,0 0,6 1.898832,0 C 35.053906,194 36,193.05021 36,191.875 l 0,-11.75 C 36,178.94979 35.053906,178 33.883268,178 z" id="rect14063" style="color:#000000;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" sodipodi:nodetypes="sssscccccscccsscccccsssss" inkscape:connector-curvature="0"/>
    </g>
    <path d="m -252.93756,649.01715 -3.56249,-0.016 c -2.51115,1.30826 -2.88681,4.57261 -2.06249,7.56248 1.08953,3.95154 3.26699,6.72334 6.18748,5.81248 4.0738,-1.27088 4.19302,-4.59783 2.93749,-8.49998 -0.66404,-2.06383 -1.89568,-3.7267 -3.49999,-4.85936 z m 9.93747,6.17186 c 0,1.75946 -0.71594,3.26127 -1.5,4.43749 l 0,0.0624 -0.1874,0.125 c 0,0 -0.50952,0.59837 -1.12499,1.18749 -0.61462,0.58922 -1.5625,1.375 -1.5625,1.375 -0.7713,0.57968 -1.1875,1.34601 -1.1875,2.18749 0,0.84434 0.53654,1.6075 1.3125,2.18749 0,0 1.5736,0.96414 2.43749,1.6875 0.86354,0.7238 1.875,1.68749 1.875,1.68749 1.16965,1.09974 1.93749,2.8523 1.93749,4.81249 0,1.68819 -0.5353,3.21907 -1.43749,4.31249 l -1.375,1.74999 8.56247,0 c 2.34128,0 4.24999,-1.89957 4.24999,-4.24999 l 0,-23.49992 c 0,-2.35042 -1.90871,-4.24999 -4.24999,-4.24999 -1.14773,-0.014 -3.64297,0.004 -3.64297,0.004 l -0.031,1.97129 -5.13194,0.57558 c 0.7509,1.3041 1.03662,2.60573 1.05596,3.63721 z m -19.99994,4.87499 0,11.24996 c 3.47287,-2.32521 9.68747,-2.37499 9.68747,-2.37499 0,0 0.027,-0.0372 0,-0.0624 -2.49155,-1.91534 -1.4375,-4.12509 -1.4375,-4.12509 -3.8524,0.3282 -5.61338,-1.10972 -8.24997,-4.68748 z m 10.12497,11.06246 c -3.46111,0.1948 -7.91464,1.6274 -7.99998,5.06249 0,2.05473 1.33766,3.91718 3.24999,4.74998 0,0 0.0688,0.0442 0.125,0.0624 l 0.0624,0 9.06247,0 c 0,0 0.0212,-0.0894 0.0624,-0.125 4.90245,-4.33881 1.20038,-6.85438 -2.99999,-9.68747 -0.0758,-0.0504 -0.1874,-0.0624 -0.1874,-0.0624 -0.43799,-0.0208 -0.88055,-0.0278 -1.37499,0 z" id="path14750" style="color:#000000;fill:#babdb6;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.5;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" sodipodi:nodetypes="ccccscscccccscccsccssscccccsccccsccccccccsccc" inkscape:connector-curvature="0"/>
  </g>
</svg>
