<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Gör samlingar av dokument</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#documents" title="Dokument">Dokument</a> » <a class="trail" href="documents.html" title="Dokument">Dokument</a> › <a class="trail" href="documents.html#print" title="Välj, sortera, skriv ut">Välj, sortera, skriv ut</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Gör samlingar av dokument</span></h1></div>
<div class="region">
<div class="contents">
<p class="p"><span class="app">Dokument</span> låter dig samla olika sorters dokument på en plats, en så kallad <span class="em">samling</span>. Om du har olika dokument som relaterar till varandra kan du gruppera dem för att göra dem lättare att hitta. Om du tar till exempel en affärsresa, där du har förberett en presentation, kan ditt bildspel, dina biljettbokningar (en PDF-fil), din budgetkalkyl, och andra hybrid-PDF/ODF-dokument grupperas som en samling.</p>
<p class="p">För att skapa eller lägg till i en samling:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Klicka på  <span class="gui">✓-knappen</span>.</p></li>
<li class="list"><p class="p">I markeringsläget, bocka för dokumenten som ska samlas ihop.</p></li>
<li class="list"><p class="p">Klicka på <span class="gui">+-knappen</span> i knappraden.</p></li>
<li class="list"><p class="p">I samlingslistan, klicka på <span class="gui">Lägg till</span> och skriv in ett namn på den nya samlingen, eller välj en befintlig samling. De markerade dokumenten läggs sedan till i samlingen.</p></li>
</ul></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Samlingar beter sig inte som mappar och deras hierarki: <span class="em">du kan inte ha samlingar inuti andra samlingar.</span></p></div></div></div></div>
<p class="p">För att ta bort en samling:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Klicka på  <span class="gui">✓-knappen</span>.</p></li>
<li class="list"><p class="p">I markeringsläget, klicka på samlingen du vill ta bort.</p></li>
<li class="list"><p class="p">Klicka på Papperskorgknappen i knappraden. Samlingen tas bort, men dokumenten kommer finnas kvar.</p></li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="documents.html#print" title="Välj, sortera, skriv ut">Välj, sortera, skriv ut</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
