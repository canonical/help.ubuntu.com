<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Snabbinställningar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 24.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Snabbinställningar</span></h1></div>
<div class="region">
<div class="contents pagewide"><p class="p">Snabbinställningsknapparna i <span class="link"><a href="shell-introduction.html.sv#systemmenu" title="Systemmeny">systemmenyn</a></span> låter dig snabbt slå av och på tillgängliga tjänster, och välja Bluetooth-enheter eller trådlösa nätverk.</p></div>
<section id="wifi"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Trådlöst</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="media media-image floatend"><div class="inner"><img src="figures/shell-exit.png" width="250" class="media media-block" alt=""></div></div>
<p class="p">Tryck på knappen <span class="gui">Trådlöst</span> för att slå på och av det trådlösa nätverket.</p>
<p class="p">Knappen visar det för närvarande anslutna trådlösa nätverket.</p>
<p class="p">Tryck på <span class="media"><span class="media media-image"><img src="figures/go-next-symbolic.svg" class="media media-inline" alt="right"></span></span> för att visa tillgängliga nätverk.</p>
<p class="p">Välj ett nätverk för att initiera en anslutning, eller välj <span class="gui">Alla nätverk</span> för att öppna inställningspanelen <span class="link"><a href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlöst</a></span>.</p>
</div></div>
</div></section><section id="wired"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Trådbundet</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">Tryck på knappen <span class="gui">Trådbundet</span> för att slå på och av trådbundet nätverk. Knappen visar information om den aktuella trådbundna nätverksanslutningen. Tryck på <span class="media"><span class="media media-image"><img src="figures/go-next-symbolic.svg" class="media media-inline" alt="right"></span></span> för att visa fler inställningar. Välj <span class="gui">Trådbundna inställningar</span> för att öppna inställningspanelen <span class="link"><a href="net-wired.html.sv" title="Trådbundna nätverk">Nätverk</a></span>.</p></div></div>
</div></section><section id="bluetooth"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Bluetooth</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">Tryck på knappen <span class="gui">Bluetooth</span> för att slå på och av bluetooth. Knappen visar namnet på den första enheten, eller antalet anslutna enheter. Tryck på <span class="media"><span class="media media-image"><img src="figures/go-next-symbolic.svg" class="media media-inline" alt="right"></span></span> för att visa parade och anslutna Bluetooth-enheter. Välj en att ansluta eller koppla från. Välj <span class="gui">Bluetoothinställningar</span> för att öppna inställningspanelen <span class="link"><a href="bluetooth.html.sv" title="Bluetooth">Bluetooth</a></span>.</p></div></div>
</div></section><section id="power"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Strömläge</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">Knappen <span class="gui">Strömläge</span> visar aktuell inställning för <span class="link"><a href="power-profile.html.sv" title="Välj en strömprofil">Strömläge</a></span>. Tryck på knappen för att växla till <span class="gui">Strömsparare</span> eller tillbaka till aktuell inställning. Tryck på <span class="media"><span class="media media-image"><img src="figures/go-next-symbolic.svg" class="media media-inline" alt="right"></span></span> för att välja från alla lägen. Välj <span class="gui">Ströminställningar</span> för att öppna inställningspanelen <span class="link"><a href="power.html.sv" title="Ström och batteri">Ström</a></span>.</p></div></div>
</div></section><section id="toggles"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Brytare</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">De andra knapparna visar aktuell status för <span class="link"><a href="display-night-light.html.sv" title="Justera färgtemperaturen för din skärm">Nattbelysning</a></span>, <span class="gui">Mörk stil</span>, <span class="link"><a href="net-wireless-airplane.html.sv" title="Stäng av trådlöst (flygplansläge)">Flygplansläge</a></span> eller belysning för <span class="gui">Tangentbord</span> om tillgängligt. Tryck på knappen för att slå på eller av.</p></div></div>
</div></section><section id="background"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Bakgrundsprogram</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">Antalet bakgrundsprogram som körs på systemet visas längst ner i systemmenyn. Klicka för att visa en lista över dessa program. Att välja ett program från listan öppnar ett fönster för det programmet och tar bort det från <span class="gui">Bakgrundsprogram</span>. Välj <span class="gui">Programinställningar</span> för att öppna inställningspanelen för <span class="gui">Program</span>.</p></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — Få GNOME att arbeta för dig, från hårdvarukontroll till sekretessinställningar.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
