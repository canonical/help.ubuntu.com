<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vad är GNOME Klassisk?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 23.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html.sv" title="Ditt skrivbord">Skrivbord</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Vad är GNOME Klassisk?</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p"><span class="em">GNOME Klassisk</span> är en funktion för användare som föredrar en mer traditionell skrivbordsupplevelse. Medan <span class="em">GNOME Klassisk</span> är baserad på moderna GNOME-teknologier så erbjuder den ett par ändringar av användargränssnittet såsom menyerna <span class="gui">Program</span> och <span class="gui">Platser</span> i systemraden och en fönsterlista längst ner på skärmen.</p>
<p class="p">Du kan använda <span class="gui">Program</span>-menyn i systemraden för att starta program.</p>
</div>
<section id="gnome-classic-window-list"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Fönsterlist</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Fönsterlisten längst ner på skärmen ger tillgång till alla dina öppna fönster och program och låter dig snabbt minimera och återställa dem.</p>
<p class="p">Översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> är tillgänglig genom att klicka på knappen på vänster sida av fönsterlisten längst ner.</p>
<p class="p">För att nå <span class="em">översiktsvyn <span class="gui">Aktiviteter</span></span> kan du också trycka på tangenten <span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span>.</p>
<p class="p">Till höger på fönsterlisten visar GNOME ett kort namn på den aktuella arbetsytan, exempelvis <span class="gui">1</span> för den första (översta) arbetsytan. Dessutom visas det totala antalet arbetsytor. För att växla mellan olika arbetsytor kan du klicka på namnet och välja arbetsytan du önskar från menyn.</p>
</div></div>
</div></section><section id="gnome-classic-switch"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Växla till och från GNOME Klassisk</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="note note-important" title="Viktigt">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m12.5 2a9.5 9.5 0 0 0-9.5 9.5 9.5 9.5 0 0 0 9.5 9.5 9.5 9.5 0 0 0 9.5-9.5 9.5 9.5 0 0 0-9.5-9.5zm0 3a1.5 1.5 0 0 1 1.5 1.5v6a1.5 1.5 0 0 1-1.5 1.5 1.5 1.5 0 0 1-1.5-1.5v-6a1.5 1.5 0 0 1 1.5-1.5zm0 10.5a1.5 1.5 0 0 1 1.5 1.5 1.5 1.5 0 0 1-1.5 1.5 1.5 1.5 0 0 1-1.5-1.5 1.5 1.5 0 0 1 1.5-1.5z"></path>
</svg><div class="inner"><div class="region"><div class="contents">
<p class="p">Du måste ha paketet <span class="sys">gnome-shell-extensions</span> installerat för att göra GNOME Klassisk tillgängligt.</p>
<p class="p"><span class="link-button link"><a href="apt:gnome-shell-extensions" title="apt:gnome-shell-extensions">Installera <span class="sys">gnome-shell-extensions</span></a></span></p>
</div></div></div>
</div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">För att växla från <span class="em">GNOME</span> till <span class="em">GNOME Klassisk</span>:</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Spara allt osparat arbete och logga sedan ut. Klicka på systemmenyn på höger sida av systemraden och välj sedan det korrekta alternativet.</p></li>
<li class="steps"><p class="p">Ett bekräftelse meddelande kommer att visas. Välj <span class="gui">Logga ut</span> för att bekräfta.</p></li>
<li class="steps"><p class="p">På inloggningsskärmen, välj ditt namn från listan.</p></li>
<li class="steps"><p class="p">Klicka på knappen <span class="media"><span class="media media-image"><img src="figures/emblem-system-symbolic.svg" class="media media-inline" alt="inställningar"></span></span> i det nedre högra hörnet.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">GNOME Klassisk</span> från listan.</p></li>
<li class="steps"><p class="p">Skriv in ditt lösenord i inmatningsrutan för lösenord.</p></li>
<li class="steps"><p class="p">Tryck <span class="key"><kbd>Retur</kbd></span>.</p></li>
</ol></div>
</div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">För att växla från <span class="em">GNOME Klassisk</span> till <span class="em">GNOME</span>:</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Spara allt osparat arbete och logga sedan ut. Klicka på systemmenyn på höger sida av systemraden, klicka på ditt namn och välj sedan det korrekta alternativet.</p></li>
<li class="steps"><p class="p">Ett bekräftelse meddelande kommer att visas. Välj <span class="gui">Logga ut</span> för att bekräfta.</p></li>
<li class="steps"><p class="p">På inloggningsskärmen, välj ditt namn från listan.</p></li>
<li class="steps"><p class="p">Klicka på alternativikonen längst ner till höger.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">GNOME</span> från listan.</p></li>
<li class="steps"><p class="p">Skriv in ditt lösenord i inmatningsrutan för lösenord.</p></li>
<li class="steps"><p class="p">Tryck <span class="key"><kbd>Retur</kbd></span>.</p></li>
</ol></div>
</div></div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-overview.html.sv" title="Ditt skrivbord">Ditt skrivbord</a><span class="desc"> — Arbeta med program, fönster och arbetsytor. Se dina möten och saker som är viktiga i systemraden.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
