<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Anslut till ett trådlöst nätverk</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 20.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a> » <a class="trail" href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlösa nätverk</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Anslut till ett trådlöst nätverk</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Om du har en dator med trådlöst nätverk kan du ansluta till ett trådlöst nätverk som är inom räckhåll för att få internetåtkomst, titta på delade filer på nätverket, och så vidare.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna <span class="gui"><a href="shell-introduction.html.sv#systemmenu" title="Systemmeny">systemmenyn</a></span> på högersidan av systemraden.</p></li>
<li class="steps"><p class="p">Välj <span class="gui"><span class="media"><span class="media media-image"><img src="figures/network-wireless-signal-excellent-symbolic.svg" height="16" width="16" class="media media-inline" alt=""></span></span> Trådlöst nätverk inte anslutet</span>. Då expanderas delen om trådlösa nätverk av menyn.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Välj nätverk</span>.</p></li>
<li class="steps">
<p class="p">Klicka på namnet på nätverket som du vill använda, klicka sedan <span class="gui">Anslut</span>.</p>
<p class="p">Om namnet på nätverket inte finns i listan, prova att klicka på <span class="gui">Mer</span> för att se om nätverket finns längre ner på listan. Om du fortfarande inte ser nätverket, kan du vara utom räckhåll för nätverket eller så är nätverket <span class="link"><a href="net-wireless-hidden.html.sv" title="Anslut till ett dolt, trådlöst nätverk">dolt</a></span>.</p>
</li>
<li class="steps">
<p class="p">Om nätverket är skyddat av ett lösenord (<span class="link"><a href="net-wireless-wepwpa.html.sv" title="Vad betyder WEP och WPA?">krypteringsnyckel</a></span>), mata in lösenordet när du blir tillfrågad och klicka på <span class="gui">Anslut</span>.</p>
<p class="p">Om du inte känner till nyckeln, så kan den finnas på undersidan av den trådlösa routern eller basstationen, eller i dess instruktionsmanual eller så kan du vara tvungen att fråga personen som administrerar det trådlösa nätverket.</p>
</li>
<li class="steps"><p class="p">Nätverksikonen kommer att ändra utseende under tiden som datorn försökt ansluta till nätverket.</p></li>
<li class="steps"><p class="p">Om anslutningen lyckas, kommer ikonen att ändras till en punkt med flera böjda streck ovanför sig (<span class="media"><span class="media media-image"><img src="figures/network-wireless-signal-excellent-symbolic.svg" height="16" width="16" class="media media-inline" alt=""></span></span>). Fler streck indikerar en starkare anslutning till nätverket. Färre streck innebär att anslutningen är svagare och kanske inte är så tillförlitlig.</p></li>
</ol></div></div></div>
<p class="p">Om anslutningen misslyckas kan du bli tillfrågad om lösenordet igen eller så berättar den bara för dig att anslutningen har kopplats ifrån. Det finns ett antal olika saker som kan ha orsakat detta. Du kan till exempel ha matat in fel lösenord, den trådlösa signalen kan vara alltför svag, eller så har din dators trådlösa kort problem. Se <span class="link"><a href="net-wireless-troubleshooting.html.sv" title="Felsökning av trådlösa nätverk">Felsökning av trådlösa nätverk</a></span> för vidare hjälp.</p>
<p class="p">En starkare anslutning till ett trådlöst nätverk betyder inte nödvändigtvis att du har en snabbare internetanslutning eller att du kommer att få snabbare hämtningstider. Den trådlösa anslutningen ansluter din dator till <span class="em">enheten som tillhandahåller internetanslutning</span> (som en router eller ett modem), men de två anslutningarna är olika, och kan därför köra på olika hastigheter.</p>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlösa nätverk</a><span class="desc"> — <span class="link"><a href="net-wireless-connect.html.sv" title="Anslut till ett trådlöst nätverk">Anslut till Wi-Fi</a></span>, <span class="link"><a href="net-wireless-hidden.html.sv" title="Anslut till ett dolt, trådlöst nätverk">dolda nätverk</a></span>, <span class="link"><a href="net-wireless-disconnecting.html.sv" title="Varför kopplar mitt trådlösa nätverk ner hela tiden?">koppla ifrån</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="net-wireless-troubleshooting.html.sv" title="Felsökning av trådlösa nätverk">Felsökning av trådlösa nätverk</a><span class="desc"> — Identifiera och fixa problem med trådlösa anslutningar.</span>
</li>
<li class="links ">
<a href="net-wrongnetwork.html.sv" title="Min dator ansluter till fel nätverk">Min dator ansluter till fel nätverk</a><span class="desc"> — Redigera dina anslutningsinställningar och ta bort det oönskade anslutningsalternativet.</span>
</li>
<li class="links ">
<a href="net-wireless-disconnecting.html.sv" title="Varför kopplar mitt trådlösa nätverk ner hela tiden?">Varför kopplar mitt trådlösa nätverk ner hela tiden?</a><span class="desc"> — Du kan ha låg signal eller så kanske nätverket inte låter dig ansluta ordentligt.</span>
</li>
</ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
