<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Dela ut dina personliga filer</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="prefs-sharing.html" title="Dela-inställningar">Dela-inställningar</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a> » <a class="trail" href="sharing.html" title="Dela">Dela</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Dela ut dina personliga filer</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan tillåta åtkomst till <span class="file">Publikt</span>-mappen i din <span class="file">Hem</span>-mapp från en annan dator på nätverket. Konfigurerar <span class="gui">Personlig fildelning</span> för att låta andra komma åt innehållet i mappen.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Du måste ha paketet <span class="app">gnome-user-share</span> installerat för att <span class="gui">Personlig fildelning</span> ska vara synligt.</p></div></div></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Dela</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Dela</span> för att öppna panelen.</p></li>
<li class="steps">
<p class="p">Om <span class="gui">Dela</span> är <span class="gui">AV</span>, slå om den till <span class="gui">PÅ</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om texten nedanför <span class="gui">Datornamn</span> låter dig redigera den, kan du <span class="link"><a href="sharing-displayname.html" title="Ställ in visningsnamnet för din dator">ändra</a></span> namnet din dator visar på nätverket.</p></div></div></div></div>
</li>
<li class="steps"><p class="p">Välj <span class="gui">Personlig fildelning</span>.</p></li>
<li class="steps">
<p class="p">Slå om <span class="gui">Personlig fildelning</span> till <span class="gui">PÅ</span>. Detta innebär att andra personer på ditt aktuella nätverk kan försöka ansluta till din dator och nå filerna i din <span class="file">Publikt</span>-mapp.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">En <span class="em">URI</span> visas genom vilken din <span class="file">Publikt</span>-mapp kan nås från andra datorer på nätverket.</p></div></div></div></div>
</li>
</ol></div></div></div>
</div>
<div id="security" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Säkerhet</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Kräva lösenord</dt>
<dd class="terms">
<p class="p">För att kräva att andra personer använder ett lösenord när de använder din <span class="file">Publikt</span>-mapp, slå om <span class="gui">Begär lösenord</span> till <span class="gui">PÅ</span>. Om du inte använder detta alternativ kan vem som helst försöka visa din <span class="file">Publikt</span>-mapp.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Detta alternativ är inaktiverat som standard, men du bör aktivera det och ställa in ett säkert lösenord.</p></div></div></div></div>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div id="networks" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Nätverk</span></h2></div>
<div class="region"><div class="contents"><p class="p">Sektionslistan <span class="gui">Nätverk</span> listar nätverken som du för närvarande är ansluten till. Använd <span class="gui">ON | OFF</span>-knappen intill respektive för att välja var dina personliga filer kan delas.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="sharing.html" title="Dela">Dela</a><span class="desc"> — <span class="link"><a href="sharing-desktop.html" title="Dela ditt skrivbord">Skrivbordsdelning</a></span>, <span class="link"><a href="files-share.html" title="Dela filer visa e-post">Dela filer via e-post</a></span>, <span class="link"><a href="sharing-media.html" title="Dela din musik, foton och videor">Mediadelning</a></span>…</span>
</li>
<li class="links ">
<a href="prefs-sharing.html" title="Dela-inställningar">Dela-inställningar</a><span class="desc"> — <span class="link"><a href="sharing-bluetooth.html" title="Styr delning över Bluetooth">Bluetooth-delning</a></span>, <span class="link"><a href="sharing-personal.html" title="Dela ut dina personliga filer">Delning av personliga filer</a></span>, <span class="link"><a href="sharing-desktop.html" title="Dela ditt skrivbord">Skärmdelning</a></span>, <span class="link"><a href="sharing-media.html" title="Dela din musik, foton och videor">Mediadelning</a></span>…</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
