�PNG

   IHDR  (  �   ��Z�   �zTXtRaw profile type exif  x�mP[!��=�<|p��Mz��(��i'F�q����Bɵ-%DE�i��g�$3NP��:hJ��2{�ϸ�qae���&Ԟ�8����.�pDF��(����!��[�h���+��|�G�NG�w/զwf{��.VV���x,�Fآm�˝���pb�7��^rY殤��  �iCCPICC profile  x�}�=H�@�_S�"�q�P����U(B�P+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�F�iV�,�鶙N&�lnU�"�D0Qf�1'I)���{�z�Y���}j�b@@$�e�ioOo��}�(+�*�9�I$~�����ό���<q�X,v����dj�S�1U�)_�z�r��Uj�uO��p^_Y�:�a$��%H���2*��U'�B��>�!�/�K!W��B������w�Var�K
'����B�@��8�ǎ�<������W��'���;����붦��;���!��+i
��~Fߔ"�@��[k�@��J� ��h���}����ۿgZ�� ��r�(˞�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:92503738-947b-4d1a-89af-b3df84e2a8e2"
   xmpMM:InstanceID="xmp.iid:6784fcd7-65bd-4965-b6c0-eb9c01861140"
   xmpMM:OriginalDocumentID="xmp.did:aac9be13-79e2-41ff-bb37-1e71a71e8464"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679601063825417"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T20:51:03+01:00"
   xmp:ModifyDate="2023:03:23T20:51:03+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:af577246-0be9-48db-ae20-af68545fcad1"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T20:51:03+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>�r'L   	pHYs  �  ��+   tIME�
*==   tEXtComment Created with GIMPW�    IDATx��}wtUו����W՞$� I Q���c��.�'v�-Ʊ��)N_�Y��&��I2��^Y�/Y�x�f�d�8�'�1�0ؔ� ��&���ӫ����c�{%@!�f�o%�{�[�>��������������qQ��h\Ep�݁@ ##����n�+t[��L&C�P8�F�RJ-xW+222rrrRRR�Xy�W;::ZZZ��x��.�:5�|!F�UPP����"��+���)))�h4�Lj��q5!++k̘1.�9�D X�lYJJ
 tww�]���]���˫���Z$9v옣��R5�px<����� 233�|�I�� �x��7�$�A�?77���U!"Z�u^o3++����{����O?�H$��x8>׸~�?''�����=�߫ƕD5jK��_s���z�������3f�p�Μ9s�SSS~�����weee�@�0���G?��OKJJ��`0����x�W�q%�0�@ p^��4͎��{ss� O����z��k������㏗�������Ԍ��ܶŋ�q������Ç��K/�}��$�0���T-xW�����������;��O>y뭷>��ϟ�������/~�v��U�V��n>8s��իW'�ɮ�����s�6�q���/��������m۞{�	&̟?�q��Ҵ��q@!�9��-��2k�,�cǎ���zꩧ�#����m���k����3oذ��GE�h4�5���7nܚ5k�������z���*�L�7nӦMx�Z�4�7�\eeeM�<������6���׳����^\\\SS�k׮s��lyN$����[!��'���_T�DʊԂ�qECJiY�a�?Q���?VUU��w���O~r��1����_����쩧�r�3��ֶgϞ�ӧ���ŋ8p���^o4=�%�b��Ǐϙ3��6e��0N�81�/���W��KKKs,�3p�]w}��_OKK����F���|�K_�RJJ�ܹs;::�
��H$�m۶�7������>|x˖-�_�ڵk[ZZ
���C�P��&�ɔ��[n�������ٲ,��=q���{,����g$��Egg'�Vk<�+�d���'���	


ؼ?~��yrrr ���d�ر�R��������>��~�>����� P\\������Zk׮���{��'�,Yr���������<���������eYΧZ�4�hQ{{{fff�֦�h���~�Ǐ��g�Ν�illliiI$�����瞫��]�d�ʕ+C������}���Ǐ�P(�X�:eL�*@nnn~~��q�y���p�.�+�Lnܸ�C)�/�7o"���u��UWW_	��Ŏ;�O�j������5j�Օ!��:=q�DWWW�闪qU��P�4M��c�U$~R����'N���ǵ�Ӹ���������ӽ^�^k�f8�Ԗ�S���i\}��+Y�qΚ�r�E�j�O� 	 � A	BBD �S  A$� ���@"
[��Y�J),"I 	���B  "�+"@� �@`��^+���O�����ꢀ���PR_�N H@����� %����@])Ӏ ���)��!��d AJ��4%"H $u�H yH$@D(��H���$DR?C�F���@��	%�wE���	H����$" I )�Ȓ�� ��K7�L@ u�� D��\!D�
���)Q��3 $ ,"�$@B�eޏᷨ��i����ҝ�D`_�=u	$ "I]٧�<�	I��P�  ��d� $	��U��yJ �'$��ʼT��|P�d�[@ $�e��Ε!� !��{U��=K�H�%�i!	=��y�,[���Ҏ�R��SA4�@[>�"XPH� ����H��+�§8�}"�O�$�� ����@�g��@���X�I��SS�{5�A�}A�δ�>��6ا�,gjV�i���WCB�ypnP
^I �(I�$߱���z@DH(��
�d���4ۋ�#i��V���7 I @h�DJ�IJ[���W��~��&�"��@ߧ-BΧ�w�?r� 	`�w�D@��z{��I )$9k�s*�K�D$�c��QD�Y\�;��):7DH���?~��J;���
 D�H�U'����-�#@�h�+��"D@��l��� �B	�RS%	^�� HR�[(I��$$�T:��@�Bo+%��y �Z>%�R �e��>S_8�I���*!��;�f����jE�d+w[��R��Geq�ms`U�V$�wd+D5/$ JeD�Μ�,)�%���!�~P`����$p����m=��W{eG����{g(��v�`�>&���ժD�	g�J�O�S�WIr�[ ��d?x�ʄp�����!(�K]3�
�$e��WR��7�zC,�K�2xmCD�#� ���Qk3 �uT����	 ��
$)�"�V�b�@H ɏ�MB��-DBr��p!�x�ņ%�{�&�H@H�.Ȭ�� ����s�g/���g-�P�8K�D�[��N�H��'m���JPv�T����g�:�p���4I8�?`˂�쳶ڋ���ζ�!���~@�s���HJ,�s���g1a�G�
�^���Ȁc=���Lp$Ǟ"�$%���e����7G��#�����Nss�����^y�&?�^�%�d�9j~����uv������Vt}��m�?�S��6)m5)�,�<uA(�ݥ�(i;	�E�$���H�i�����I�3nu���������>&��p؆�2Z���'D�ñF쥻�lx�#�+[}���i�,�}��Ǘֻ����]�{�{��V:m��>!��\����g�H}.ԹzG� �s��9N+J؏�6P��|��)SN��	Ѷ��P�m�e
��2�D�	a����mx3�p\>B��,�i�M�cI�$��c5��,�x�#ɎM��'!
�]g���@�/޶Ӕ[j)M�L$�@Xʓ KJ)�2e"��&���G#�Ƥ!����U��0	B ��!��,O2�7�.+�R��t U�A8��c��Y�S4�WE�]����(�� ��5)�� Q�$i�)�)Ɋ��m�}=�1�Ӓ��4�O�`!�o��qI�M&<ш�$����
��Uu}��1���� P8�Z���pr�C�O&@�)-�L�[�͑ݡ������oK�S-�����<^O�ǟ��%!���8	���:`��wⷤ|aLpv��{�^{|�H�	J�E�tDk"���bhh|j$�"�
�%�$�L7�����;�����NV�Ҏ�	�Cqhoh I	�;@D$����fGstw{d�i%�a���?��'-3	q� T�"o������y�;T�&�N�QE�﯂Ty%la�i�I4����ן�yWC�S-~1��a�pj4��R�Z��I7�M
 v	�P�J�`�QmZ"�&3�$�,JD�=[C�zm^jh��O#�Dz� O�� �ݻ�Vs���>��/t6��H"���LF��-�X�6/54�2�OA4�u�"��T��(Hp^ )Cզ�D"T����J: �dYVҌ6�|���R��q,���F������鐢��D�d|�ʪB@	(�<� B�-L3i�4E�wF�jSC�fg25'�J Ke��I|��Po�:�<vZJ��,)������A�S��1��'e2%-�v^������N v�HHN�DU� 8'��%e2a��{v&ͨ~�˞�y�q{� P�ܑa\Щ�8-;���&I������X�cȮ3�9E�N��Ÿ�K9�����;���p]�cY�@<5H�5@�S�`gq�����0�H��ҊZ�]�#�e�~��K�<*ƲF�Q^ʱ4.��9���~��@�YI/�XD�r%=�D��w�\v��N�r��E�D�ʴ	,I��f(q"�hA1��p��ĥK�B�r���)~u,˲|�d<f�tT'I��L����{v�E{\��$�;~DJ�$��r�q�i?=��x)�Ҹ���Bߣ²�!�N]��P�n�L�$���	$ �A �� ����m����bf{4�2x!�0c�w��Y�i��q�H��!��K8���L�A�$�$�Y�g���8ɛٯ$"
'�%����1^�o/�XC����å�p�xZ<
G�q���%�6%�$����Q�q�Vو��A2u_ʱ4�X���3\ʱ��eX(,I���)�`f6�?t�	�4����sAA�	4]Qci\T#sD^����K?�#}�[�1'�p(Y��PtIh3I����26��`�O=OVV�aD�����8�yI�ϫ��@fff(�c� �Ҹ��nD��=�wΜw����D"qF��!��(=�[�a�kZ�� ��\����,�I+�l�\H�������v_s�5��r��ٳ�M�fFSSS2����0��5MsΜ9+W�LII9x�`jj�iD��2�T!DAA��������� �5�m ��cq�;�����:uJ1��x���+uD���o6#�p��QB2M��`J2���{���`�ܹ999n���?���3f̢E�&N���޾cǎ�G��}���б��f͚={v<���BL�4)z��C�UVV:=�?����ym�����K��bʔ)���������v.i`,!Daa���_�s�Δ��׻hѢ���������!��wAGI0Q�p4W�T���^�G �	�i��eɒ%iiiܲeKkk�	���6m���A�o������:���������=z4"677���ѣGggg��坫�� ci\l�7��͛��Ҳf͚�����g���C>� ���/_�<�����cǎ���/[�l #n�sF ���Z;�մ9�������"y���!77��?ܵk׬Y��ϟ�v�������,**�뮻�mr=��l����ҲiӦ��v���7�3f��!��q�/##���áP(G�ь���!x3f� ��7vvv�<������\�t����:4�sj]��L؄݊a[qn��(�nD�h}Qa�fZZZEEEMM����>�`���cƌ1MshQ�s��|����r�4w��y�ȑ���S�Nmݺ5��Z������~U�aEEE�a���͜9sƌ�@ ����X���� �Ν;��ꈨ��������t���;B/�9ף����B�W�W�����'N����ǎ�x<^�w`_yhO���G��H$���b�x<�������q����s�-�x��I�&M�4�Q�+V�x饗F�<�����O��4M��;�S� �O�Ǐ�(�� B7�}�H���~�3f�X�|y[[۹�����[o���{�ޢ�"���oNKKkoo��7�
��e� ���[�A����5??�w.###55���u�O�
vo�ʧ�����n5|ًD"[�l���˖-��7onkk�v���cǎ@yy��%K���,XPQQ��555:z�q6���?~�����Q��ӧ���8p`��"�F�Npڹ�(�k>��`4]]]cƌimm�R~��ǻv�R&��ѣG����B�~�ah5�n�;== <;�9%QJJJ �����4FD�l<y��s�U]]���}��7<x�رcn���������?@=~���4��ե�ۆJ��N%��4::�"����^?����痕��}ۡPh�Ν�:]� c%����o�H��������������?NOO?~����L-x�R�sE�L�L$��l�i�a����>����{ҤI3f̰,���iÆ�g�w�������/��.��!
�DɅ�ɤk����2�1�B���.�+���eY�H��Mm�4�\c9�˲&O�<��}��}��G��<���"�+O�0���Գ?�,�\9�R�~��y�r&���s��D�H$�p��:m����)I�p!���HB
��M���Q�V\�{��bY� ��!������w�a�ci\TS�\Ƌi����t����r&I����:��T'������i~N�Nk�z&�HQ*�.�X#��/\ʱ�|��	/���6��ux`7��~�HC[��o��$�r,�+\���.�X}t^o�l�ds>��{$�PJ�a���������R��qQC,����K9����s�;�	��c*[�����!�*�a�����ci\T�74]DD:.�X����凂�T�
�P'	�M$J.�i��L�̺w)�Ҹ�doȫ��M��� @��(�5,H"pJ �dGXp�ϑ��\���K�bۜLj2����I5/�X���.Q08�io���
�H�5!�
1�� g�c8�-�T4�R��q�U/��K�?��%�W9R1�K0��y	�d+ho��]D(A����_���+C�\ʱ4.��W���W�X��.R	d�@� ��WnMi�Q�;��oNO�O�~*�"�w�;\��ݥ`�%��V��ACc�*O՞��0�#J��1�-�b�ӏLCc$OY���fjS���;r.��o��##}�1 ɖ1 ��/�w_$hSSCcD�S2�g��1��M�P��y Z�44F��D ¦n';O��@2�-[���<���\!2��r6.�O�t���#(w.��0���
hh\.p��i�#���t^DC1<�U���P��GB�<���s:Hj�Ӹ��&�h4:�C�[q!���\I�N@���[�`����!|>߹x44�P��n}�v��~<�D"7�X���8� 	%	��r)�1Bd؛C�0���4�ǣ����!���w�ݑH$�U�!��� �@w�9@�J�Z� (���������t�q�OX�����g��$��A$ni"���#$�Ү��0x�^-u�>���ZI�Heh�vB& � �\�GH���"E�z����t-u�J�����bu�/لc���w_��A ��>!DJJ��:�O1�~�P;�(&i�@ �w�� � ���L���Գ��+�}�VɆ�Xոb�w�$�m�� �B&�f�I�
�m�(Aw�݃�>Ǵ���7��-u9˲����MC��Z�~��i�� х�2���]T�	�{���%�[����2�"8���O].����L�Z�4�@����gPv�3�v����̓����l���`K�����������F��kh\b��T�E�g�6Ņ"�c�F�<�hgo"JT=�'x�MO��� ����@ Z�f����;ؙ�L*�  ��D���.�~�T�*!�E�W2���.�Zϲc��N�Ѹr�>�`��]�L_��AD���+�n���2ȋ8�M̽��l�4��;2�54F����'@�証&U�'U�9�D�����7��q���n`������/��o;55u �.t�BC�"��ch�%@��+�(��b��sd3t�	��;��������p8'''77�wH��p8|.�6�H跮q%��|�5�� ���.�����|;��w��
x����@�����n��֝;w�[��O��x~�ӟ��?��۷o?[�<����F�0���������Ś��������=�;���ɓ'��?��G?�Q<���~֯�khO@�]�;A��H��� �f��"pn�_#����y���s 466:ǥ�����Ǐ�'�n��M��nH��z<�0���e˖�3���tuu���[�=��رc�͛�u�ֺ�: HII),,DD��7a��]4�qQ�#  �!�}; �Mx��$��7�s�ν뮻zzz���?�_�~	��eY�>���w�}�w�^��СCǏ?[���y�#._�������}��g��xAAASSS"��2e�O<���ʂWWW���~7������_�su������R�������J[qvԁ�y:O��v�϶B].��ߞ���f͚��z�Ĕ����^z���d��ٷ�z������\�~O1m�4!�_��׷�~�9>~��믿��v/^�8##���6M3//o���^����q���|�Y�f���̘1���VWW�߿�?
�]w]^^^CC�eY�����?�    IDAT6l�F���\VV6~�x���'���8q�u�]w�С�>���&L�0���۷�����1��M�`�iQ�^[��ݦ��;�`nn��ɓ#�țo��R�C�P{{{,�x<��o���Ϙ1#--팤��ID����v�|�����������H$RTT4g� �7o^qq�֭[����eff����G����B_�����222���S�~��_�ڵ����[�Z�h�"�y<�S�Nm߾��Y�f=��}O�����>����ٿww�m��v�M7�߿_O�Ϛ�G@.@a	�%�E��\5RPq�!7�8�R\\�r�:����G���~��G�ю�>R__��Ԕ�����w���+�CD���ZFF���_��o|�+_��'�|����WVV����}ꩧ�~��w�y�4�H$�_��ԩSn���'�X�b�믿�{�n HKK��_��nݺŋ?��#.ܳgϢE��.]�}���^zi���_��Wθ�����q��^{mϞ=(+++((���ӦM;x�`uu����1�ǻ� @r~���RY�dI�E���"�3,�;��;�i���@ 0��������o�v�ڙ3g�|�ͳg���W������4�eq`���#--mŊcǎ-,,d=�d۶m�D"_��333�nwII���w�ݿKK�w�qF)F�'�,kÆ,�0aBKKKaa����A%�i|��<1�V��|h�A i�	BӔA�ZZZ `���令��fff&�ɳc7
D�x<^[[��+�|�߬��;vl^^�x������f͚U]]���������!".Yr�\����Μ9�n۶���aٲes��B�Ɖ�gK�;@�㗒@" HU���@�FB��۝����Hd����Ǐ?��3u�����}�����-{���o,..>x�`wwwQQQ^^^gggGGG0�I�&mڴ)�O�4)�޽{Æ���Vȷ�zkSSS~~~^^�c'sPg���g�0o۶m�ʕ�G������������z�� ��?��cJDD��RR�S�#.x�pxÆ+W�\�z������ƾ�$�())��{�hݺug�А�������|��)))�a$��������ѣ�i�ر�;�X�|���������'O>����w_gg�#96n�x�5�,\��׿�uwww0���t.[JYSSS__��c����}O��+++�.]�����{����Ϫ�1�-�ʋV�B�|(���DR�5�É筅;��/Ʊ������Ң�������6'
�p��իW�=z�Ν����قgY?φi�����޻w�����������Ν;��������ȑ#;w�<x���Çkjj<�u��W^y���v߾}����d�ȑ#UUU�p��s�Γ'O�b�ݻw���UUUm޼����4�7�|ӹ���F>aee������ښ����N ���jllܶm�Ν;�u�W#���y��ݱ�Q D��/�v3<n�L��*DD`Z2����}�B��]�����i�j�3
!�N����|'77�����ѣ'N�p�\%%%���������É��|OO�y��@zz:3mTTT��?�î]���_�E��~����uީ(���9A h�T��G.���&o�IT���
g�IK)����o��o�V��;w��ٳgϞ�?���W_moo?�lR�x<~Y���唔�H$2g����ꫯj�Ӹ s�P (8=PI����w����i���ج�������_�ZZZ������C�����K�b��eq�����˖-|��g�v�ƅ�W�� ?���!H��<��ic@H`�eʤi��c{O�����{�|��d2
�����fjf#�Hfn'޼���b�M�}D�L�FÇ^#3�h�Ӹ��%yȦ�T%�$��uB��j;R� 2g�eY===Co���qe� s������T�. �B�������A����s��V�-H	� $$A$	� ����!�6S����r�`�楔�DB[�W9H�v$�۽BoA���$0�-�ߎp��4�P(��z���\�'�L&��x<�L꨽�U/w�`F#R�SX� 	I��(S�U_<g\�08��'��)��"��p�za I��@����P"�  �C��.�劆����C_$XĈ	���$'�K��������S�+�B"�<ш@���W'	�@Os�kh׸��$���d�)Ҧ~`O�z��jhh��d���8�B: � �� A�P������ʳې�ѷ ���B��z։YCC�r�؎���R�h�v(� @ IhI�Ʀ��ؚ*g� @`�v6,�( �9�I��m�#��*#�$P�0x�ApI�HtN����Cp�9!qt .�f�X�@�����0�hhh��D@ �݀U�<A ܫ�H%m��y����!@�(���mw�SJŰ���1|�cM'a�D1`�h��&ٹ,����<��?!T�BA�$���nBN/�y�v��?�;;S	��0%JNl�i�#��j���_Q� D$ B�,��ih���C��1��㶃�D��E����[��i�W*�M�>�$�;Q�?%I���dK(6��	��W����T���v����o644�~��>�o�'N�8�W999�a�K���O2[��իC���w�����tn�и �w�@w"�  ��;$DaW�^�D�DjB�Q�eđ#GfϞ��x  ???33���y۶mG�ݱc��Ç���m��v����Q0t�݉D�>hnn޼ysSS��@۽CE��$ݽ1KN�$ H���A\��,\�0677ϛ7��?N&���ϟ<yr(�������把�)S��=���Y��4�ŋ�p����k׮���������_|������-Z4nܸS�N���k���>��s��ܔ)SZZZ���_}�����+V�|�w�}w׮]��LcxF&{r(z:b��$$������D(	���M\iii	��cƌ���3gά���R�ر�g�ٿ�]w�������Ə���������җ�t���M�6��⋯���'N���_��СC��{o_aӦMO?�t2���曅��~{JJʯ��cǎM�81<��o���k���jժ��4=w4���q=$!1eB��t�T�E�H��ӗ�X���S�N��b����n./Z�hҤI���l�;v�����������[��5q�ĩS�~�[�r2��l�ҥ��������^x����ݻw_s�5999ӦM��{ `ҤIڇ]C�tK� �� � $�"���2��w^s�	��]��z��cǎ'�|Ҳ���* ���������s�UWW�u�]}#:�dRJ��(���bo���_��3N;a�~��矯���5k"
!�JW,;|��3�<
�������g�@B6�
 Y	Jt'=IHH @$@D$D�˝$����DfϞ}��q >�������(55�ߟX�UPP�v�8p���������l�u>�/55U�KJJ|>_<���]�jUvv�����[�.\��������ϑ�g��T皘s�@p�(� �ҊY�E$�Ef$��^����o].Wee�i�===�����z��媫�;x�`JJ
 :t�U��ݻ���o�ᆢ����~;
}�������뛛�Y�v�ؑ���|��p8|���������q���z�>����nڴi߾}+W�����6s���cp�	�x4A 
D�Ue����!��e�]n0�$e�5R]�>��xW�����������$���`��DJ�c�Kp+f@)U���I�A���f��>�)���̜>}zWWג%K�}�]-u#ih�J����J�?@"�	+�0M�L�_�����7lذg�=W4.�ׄLhK܄T� 	�w���HJˢτ��B������sC�EW�#f0��A���Lc�����9��"9͖��A��~���544���{�<�3�P)>�����������1l�c���]�uH a� �Q���T�
+=D��q��+�Tu��R9}uV��ư|<�lD�޾S��H`q��qY5͘��0U^��I (&[)��U���������S�$!� ���Ȧb# ���/j�����lsW�I���#{���������gW��@��|�)� �"H*�[M3��1B�G�mHDo�
���T	c �����HY��� �[v	ٟ�@� �T��Z�ih���C  {�N���@�$S����y��(�@pJ4![�$Qe��*ӻ���������
����R��r�ȴ+��k\!^"���D/�x#���ezY�����x '�I�0�?^ZZ�m�6����JJJ6nܨ߹ƕad���RN?J�A$;�HHI��˛6mZ2�|���ɤ��A��ӧ�<y���%;;���E"���V�4����(==���}ҤI,8|�pSSSfff ���---�D�9yzzzVV�eY�N�2M3?? �~(J&�����e544h���0���� �H��:��I��2��ej�������ӧWUUE�Q.7n��ٳw�ڵr��������5k�TUU�{�999�pxݺu��Ņ���7o����~AA������}�?sss��"���۾}�[o���o}���ɲ�����'OJ)KKK���?�رCO��ɝ]�蚐�̩�Y ��$�D��8�E��r�����'��U�V-\�0�L:t�����?��O�h�ȑ#{�������˫�����8v�ؚ5kN�:������"��ѣG���#��6m�Ν;-�B�e˖Y����/�ݻ�������k֭[�~���ӧ?~�O��������?�3G�_�eLx�X
�`�#;5��8���dI@&b�l�F����ƍ�Ν������;edd�|�͆a;�G{zz����v/[�������z�^��u�\�w��㍍�����`в����H$r���X,�H$����͛����0A\�� HB%��@����v�;���M]a��d2YYY�o߾��\v�F�����������n���VXX8cƌ�k׮[�.��R�H$2f�Dt�\���h	���!�u�\|PCc���  $
R�T �N" �ܱ�rF�g͚5w����֔��`0�s������+W�x㍡Phܸq+V��2e�٭�������/_~�ȑ`0�bŊ��|���^ee��ի1''g�Ν���\�ҥK���^z饼�����?�yOOϣ�>z�ȑ��{Osj�O�@�( �U���q� ��i�ű$��Dqh�^>/�2ahss�u����;;;��ۉ������^JYUU�o߾��ή����zVk�P�����v3�4"���TUU����tvv>|���;v�>�R����<y2���ᆆ�m666677'���ƶ�6�4���Xg���www뉥}���x� �x o��3P;��SJ3�;�e�iQ��j[��&i��c0L҆+%�5N�@BqA�>��Z#"v�N����
�5@�NH:�
*i��n&�eOCcx.�ڥC�	m	I����;�×=D 0P�KǁM%c�G5RoTCCc����'�Ԉ��B��*H���44F��cn#�_ըR��� B$r�"�%ԥ�#dm�:I�d��� �/͍�AH��ô2""
D!�����*`9q���xÔ�^!2��@@@B�>&L�\�y�54FB��v� 
T���\�g����u��B�
���& ��؉,L2��u���0��x\eg��Rok.�,1��w��t������ET4��N�@�nK��1�'A�*�MM����'�$�$� "	mhjh����	���>�lx"�FAv/�a����d���<.�ED�$z�Z�44�#w*� �PF&�tI(T�W�$	��P�������|ɒ%���G�}��W�#�4ʹ��+Vl۶�����O�:�_�ƕjj�7�KͅJ�D�� \8�I�=�2eʔ{�g͚5]]]����drɒ%�G�~��M�lll��bMMM�x\�]�+Y���G:�do�"�T�&T��e��c�6778p������������?�4͍7���̜9��ѣ,x.�x<&Lhkk{��w���ǌ�d��˕H$�z뭮�.D7n����v�ܹ}��k��F�cǎ���y���ر���KO��u�UJR@@ ���I}�3W<XZZ�裏������twwWWWWUU�_�>�H477WVV^{�-��ӧ���o޼y�ر�V�
�_��[ZZ�9�jժ��T�i���������C���E"�U�V����[^^�	�5.Vp� ��tE8�I\v��.[P/'���~�_���Gy��_�:�H�B�������#G�������"���ݻkjj����c�"��￿u��'N8�<z�hOO���Eıc����
!Ǝ;nܸ�'O�����1N?�r<N��Vx��#$�L#m��+QCCÚ5k~��_���Ϝ9��������J&�Ǐ?CM1�_JJ�i�g��	!V�Z�`��S�N566
!�����8q�ԩS���4I��E�x�vD�,cR����j�EW�6BnnniiiJJ�aR�P(�H$����^oqq�eY���#�~�srr&M��������=OYY١C����N�{�Θ1#--���N1y��ѣG@ff�̙3].���9s&�CPy`w>7��i��99ű�7��
��ߞ���H$jjj��ߟ��z�w>��o���M7���SO�b���: 0M��?���g7o���#�tvv�5�?J$۷o��,Y��x�`CCC0ܲe�����,Y������������n;p�@ ��;^~��p8�'�Ɛ�T:���? B-�B&A �  $K�,��v�uUڦ�����?����N����65�]�B�@t��S's�	$I �Tτ��sE1f̘p8\VV���~vc�K��@"�A y�\p�
!�������zy5�'N\�hQCC�K/�t^�{��\A@���1��$�hK�]��W3��i�6lذa�~��_��RXaS�IUm�,�P���9̩��1|sS)1�~����Y�m�i554FB�B t�@Q�! H !�����P-Z�44���%��Aؔ�U�,��ֹ�:��6$�P�	A*3S�1Im��b=-v#di � �m�?"�w���MݦKCcض&��\��jW��jG��(�"�$R\,��z\�N4
H�qr+f���P7�����is?� eG�P
� DDBD�U%h���Y�ӐjHJ�� %!G`�R�����z�^��5�D"��4dqC2l�����[��BG?���f%������a  �	X��q�4G7I�N�ᮡ12n�sk.�d�qLS�nߡ�>���1d�c=���Aڤ+��)�?)T�@�:OCcDdO�g !GRx玄D ��`�?�:SSCc�b'�$�H`�U��WP��hS�� � g�  (���� -U��! '����1�g�>��H��tv�[t�s��xv/J�I��{
����ZNQۢ�654FH�q9,+:;����'�>� Ԧ��ƈ�ݴUs{�����-���^���1�`p�4W��c�f�vX ��(HCc$T! ��	��>��!��O):\�Dt�ݨ�]����M)���/ W��Ŀ��f~~�~������=P^^��ɓ��и8&8L  qjp��b�B	@$?#c'N\�x��#��Tt S�2�Ipq��ߕ���rˬY�<�o�QYYYRRr�}�!�֭[ׯ_�bŊk��&�Lfgg��G?Z�`�����M��x�.���������� ����g�Y�t�iӼ^�/��[1k\��3W?�8S8��Lw�;�WT��3ƍ��3����?��c���{���O>��'N�<y�o~��������D�k׮͛7���~��۶mkllt\G>���noo߰aCcc���{=A4F޿�2 ��JD�L5�����
 ��P@�q�����ttttvv677������n۶�4ͣG�fdd���577�J��    IDAT!��("���,Z�(�|�@ �g���16	���TE����� H i����`YVFF9����v�\}�&�ɴ�4�Aljj�c�=��'����MMMNt���n���T�I��C��*{��B�@ B��?���!\!lG^�������dܸq�5k��ٳ�/_�F��۷w�������� >\ZZ:w�����gdd�|���M�>=++�9g"�@�ٳgϘ1�C����EEE���~���;�3g ���<��Cn�;--��.((��GcH"G�vWI�R �b<��v�  I ���F:_�fjj���mBL�:uʔ)�&MZ�~��'�͛'������H$���1c�L�:[ZZ�m����0g�n�������]w�u>������ѣ�6�H444̞=��r=zt�޽���~��ԩuuu���������iii�`�СC|'N������H�A<?/�3Dt!� o��p�� �w  I+aR<�;�߮�V�h���������DTPP�}�?�!�$o�����bN�v�hp#��,m����c�A��~ ���KKK����x<����w��@ p�7��{��w��i\	�	���e�"sR1��%�����\������z زeK{{�auuu�G�~���8�_�ƕ%z@��cIU����b2�+[gtttlٲ���i��������Uk\AbG����V�|T��2�y�yc:AYCcX �D����r��W@]��1|���A���Ih��R�,R$��	��j<R�EDFo��
��jV���!i�#�a�}�H�����L��4U���:���^��&@�(�Z@@�$Ο�j��44����\�v#f66% �D�$M�}�544�om"q+fp� $!I��	^��MCc��G*O��S����4	Hp	: I-w#dp�L��"m�j�e!����<�.���Ȩ=�jD@@ Pi;P�dHDP"�P�K444���SH	U�.PD�R9|�P3Ikh���)���hgc��M;������jjh����)`�B��!��'��&_��rw�u׍;��.������f�;v�3�����IYYY�Ǉ�������gffΝ;7%%e�5�n��|z�i��� �P !JA�j��T?��{]vuW^^�x�b�����w�}�a���YYYcǎ���>�'S�L��z�����@�������M!�]wݥ��4����v�;BՅ�$�  	�<ӗ=��u����/==���kΜ9�nkk;r�Hnnnkk���Ø2eʉ'����L���������Y��w�ގ�>����L�[[[8��'N��r�rss{zz������S�RSS���O�8���ɓ'��'�P�5*"���vvv�߿?�ggg3�{JJ
"�3���8�����z'L��r��ػw���)++��|���---�F��ai�$��@�`�IP	� 6�4^�V�,H�`+***++`ڴiYYY7�|�m��f�̙3W�XQPPp���\.�S�L��Ξ3g΃>�(+&���ͽ���gϞ ˗/���;�����~�7���/_� &L��dɒ`0XRRRPP�z��I�&�m��v뭷fdd�{�s����ȸ��&N�XVV�x	999���_���@ZZڷ���n�)
!>��ϕ��~�_HOO�s���h�ҒÛI��Ub�?� �y���G��6m�eY�@`���D�v��Q�F�B����{��7�x����رc7m���Ԥ����{/77����?�pvvvCC ������;�F�JOO///߶m��-[��:uj��ů���C=���5a���'O�_�~ԨQ���S�N����Rn޼yǎ�htڴi�x�0�5k�H)�O�ND[�n���KKK{���ǌ���Q__�����MMM���˖-{�����3���4]�g��d>12ؕCn�B��t(_��E3B\.H)��ݻlٲ����a��GG���""D���ܵkתU�^~�e�rs�\��������4M��6??��;�<u���w����D��ى��P������ //��?7n�������=��N��!���B�P"�`v3!���˳��������˲L�$�@ `F04Ms�֭���zJ~f��I'+Q�����ޥ�Ef��2�����5jTEEEMMK��ɓ�}��={�0�a^^�̙3���{�u�!"O����s�[�n���D����v��{�#G�X�u�p�h���n���n����~֬Y�Xl�ƍǏ�㰥�e̘1YYY�@��o�.]�q�����p8|Ɨ���:::����~��w�y'
����o dff���������d�t�<Uj.� �$�D�	�"Ӵ�Ҕ$/�F^<߳gO~~>�����[���c��X��{��z뭻v�z��W+**���92s��Q�F555=�����{o_n�������Gy��k��≈���7o޼�>��4�cǎM�6���6mZ��?v�Xkk룏>�����@ �<x�K_��<p���i�o�������#��\����ggg��`���;����'N��W���_���<aY6�_HuR]� HJS��Ȣ�%בN���ڦ�����655�e��榥��b�D"��ٙ����������:::��yyy�������x"����H&�l�����|�h4��:::F��F{zz�^oFFFkk+�F777��q�۝���v�c�X$���{��:�+O��e����	��DR�ږ%��ͮ�r�D�[G�D���<T���<�_211S�]�����,�Z��&Aj��Ď����Ι�o���E�yD�7�����;[cyyyll�V�5�J�R�T������ȈQ�ƈK�$�"c莌���͙�a8::Z.�����;w�hll����q��,--����������|�����Tm-�G@�/O��@ ��L	3�� #hi'5��0���X>�#�����x"���l���NX�w{@j�L��9���x�#�;s�@L��@�) :-�hT���2%���$Ir�$����6��'m�L���	�1h��!	ٔi��H�-�6g�|'rz���;d<�$I;m����f����;65��vnm��PQ�$F�604}t�L�5��l�v7J��}�9;��ֺÇ�)�oEQԡ��� �&h��JtS�`G2CZ�ޡ�����(ߌ�;���g� 9]��93�DW۱��j�:5ys��kN�F��ӎ)S��mX��oA�\��T�uJqo��)�o �q�j�:����d&IҪ>�E�"�$&��^R�׳��9���#���]���z�

aZ��"(�F��>���Q��\��r�%�o0�5�����-ywOL��wLlk[ciJ�M������r�{9}S��^�w9s���!!�Oc mKv%�@���	�v{ee%����T��z��m�nJ[9"��H�Ѥi���(��$l�� ��$I����0̓�s��S�$�Z���݆�g�-&p���P��Y��31=���5�Z///
�j��a�y9}����f��܎g�x �1;�Y	!kf�m���,[~hS5�a�\����{9=Ў�!�b���N�D;�1p�'M
)E���N��.a�{�_EQQJ)�~���`r3�<�K?�!� A� )$Ƅ�5� �\�3�Q��Fr9c��Mm� ���'(D���)�b=? ;&�q$�Ġ��D�An�ӶMM�c��N@@$��] �i����nxI�i�9�ӽ9τl�.�@H�آ�akb�9�];}ѝV� 2�� Y�m1,H��)�Px�V���ZW@!���^��)s�i��O�	�"���a1+[��Ob�)���5�O$��( L �Ȧϴ�b����JN9턪3�T����Cٔ2Թ��)�r�X 4I�� ���ßx�3o��SN��: $ "�*B��֎iv͎�U��ZN9턵)Bڪ2��l7i d2�'��l�SN;��DD�	m_M 0?3"KF��>^N9�g���\M�L'w2��m޴6N_�l9�M;ӄ��t7`��)!k`�A�E�9�mB�v�ĩ3!`ad����tɓ5s�i�v�x�r��}���#���Ъ��r�i{�Nl8��İ���0 dAq3���2�)����yh�73�U���V���f�a^�SN;`jl,�i��;�RP�L
��xzN9�-γ�NL��-�e?2�����9���ؚ��P��*d��Y��Ǧ�J��r�i�|'n�L	6A��ŌB4�ʓ�r�i'�<cm�����{b*��ڙ�D<x�`��~��ĦT�T&&&FFF�hqq����+++��|��@@��1 ��9؁� ���9s��^���|�嗯_��3��I)599���}opp0 �Z�[�z��ϝ;��`�Z���� !Wt."Hi9�U��j������+��ax�С�_~yvv��C����G����?����	�`hh襗^�Z���}����JA]^������W�ު,�˃��/�����"���OOO��׿���S�Px��\�)ógώ����uWP�mwcE� ��A85
0� wR(
���p��a?�7��B-Wwae�a�,xp������:88899�l6��h-�v��ES_�(5�DI$c\��@6�M�f��B���: x�g�?n~n6��������=�����4�p��*����� ����z(iN;A�VkiiiK���Q��4Y�LiW�纷3��`�|�V���(��?!]8��m�b����鯬���U��`��h��bRW̼<�[MԌ�hjj�رcJ�_�����j��;,>�o�=�L~O
�5����م������x�N�E+  �ԙ�M���P��?���o��?��O�R/���O< /������/�˅����FsA��ٺ�ze���C�m̖ssSSS�V+灯�� �v$��"Ȅ����6ձ6u��잘9��7�x��ŋ"r�ҥj����``` ߆�����������쭷���O9=��`�D��:<��-tE�s�lI �����[p{k�m�ݾv�Z�P�p����̉'���s�|'�C������}}}�R� TQ��������t�R��}툰7�x�wzP���$!Ht�Ҫ��e�h�0"�ٳ���wjj*ߌM�T*8p```��VVV�^�Z���e�:R@���~D"I03�ġ�J@�-�)� ��i�� B�n�ʷ�Cj�Z�.]��������0<t)�@�J�����:�CF9�3�'h8�x.�fH�����H��,(����i9>2�����sn���ȭ�j�SN(< 	\�MF;�4�4�Д��L�SN;�u�&f>� �u}cfr��9���<�#B@4�K�v{P�զ-KGɻ���NZ�d���(���<1IX��r�>Y�2 M�	� f<��q���Q#Z�U
����p"��
���$idq-�EqMs$A��)�m3��.Q�ƮB��HV[I�9I�|��r�i[��	@A5Р�8j$�D�Ңt٩ :��N{(9��w�_�HP�T��]�j �fp��M�O��0ID�I�H�m�J���������(Vưw/�� �A>��XQv��Z�&7���i�rK��H�V��4���س*�VQ����$f�Mh-I��ސ����P7�#b����p�HQ�`��r����q�ѓ�{ =g�z�����w��s���m��B/����X�w�#"B�BX��q9.���,}��]@gBb�%i&�z��Q�4�
 "#�f�[�QP¡c��[�~�&����?�,~Ѻ�&��/�U8�{��a%_�-�*a�^��2�gi�ގ�	 j��X+i�0�0��sIҦ&�AX������/U�Ɵ���9�y
Җ�*DR�!Uҍ���A�=gi�S���߾)��~��Akڵ��'�f/ "�@����g��1�f,��5eKݎT��=��ǁr��1
��U&_��p�n�Y;���ގq_e����[a\;HĢ+�H� ,�bF1�h�ڕ�I�����ܗ��MW�ҁg;2q�=	����m(�����toe��*��a��i��K'�w!�p�P��З���v=�9;�}���\�}Y�W�]g�:��b	 @llK;0�gg��cW�
*���ŗ��
c�Qy`�n���r}y�N`Ϟ�O��3q<���̿�+m)��*tl4Vwcel�O
�}� �f��|m���"L��׿|�о˦�B��ph"j����a����}_8V�S�S�q�yJ7VppRV�wʪ���3��bv]\7��#6^^g��@��y3ҫ��Y܅Y6d���j�'5����b��Zc�~w��w x��;i߀pߠ�E2W�GF�Z$�W�V���~*���������Gʯ_n^_H6e�pd�=���xc�wz;��}�R�C���W�(�������@+�۫z�� �Ȯp���k܁@��Z;_vDd �)��Aui6�d�0N��7@�;Rx���"�Zڊ��e4X���;�5�2��v*b�Ppf�GK?x��̡��}��2�}��w@��=\:: �w��ٽEd�[|�`�Y��ॆ��di�P��)�Pe�^�VƺB�jm9s���#�b����>T|n���x���9Y1�7/+�|a��;V��bv��W-� c����B��P�w�b0	\z��( �"�@b�u$�0(c���O�^�S3�ݡ�a�ϼs%z�JtbO��å�|�Xnj�է4C!�vQ"_����զ}�R�#=�\@�UP-Ё����|�-#��fW�`����xO�j�R-b+�;����^*�X)�g�᪲��i�7���6���_�����O�?ռ2w_�G������OCy���w��צ����x�O�/\�n��X��%���<�'��c�b�Ͷx��_�,k �SwVu��Y�f,s5=TUca1���,�`�G�B�E��ЦQ�H��1�e��,�0���\J����ҏ�(DXi�b�S|سGVot�u�H   ���n�͝:$`4�q�#BP��7������Á?}�:kcMmL_�_�/<7Q�\�����B �X~u�9W��O���m-C�<k_��H��OU���O[�?}�X��'�v��_�o�g*KM)��~�a��Rrr<|�p)N��L� 80<?Yb�B���ue.�~�����z��'����s���N�XZ����{�tϠR'�ʕ;�ɽ�ߜ�<�����ۥ�B}��W�C���~usIg�с����+���:!��S�_|���,1C!�7.G�V�oP��e}z_���E�/�z�ye.�?�t� � ߹M��{�b '��Ä/+��p����Q�=X��aO�"W�`���tLD�١����I&�x��X������R] �>Vy�D
���۵;��c�-��_��HBW����p�|x$H�[�����U�ÓeoYOݎ��Y�����7ЮJ�뭙���*����?q�85�~�J���ˁ�b��(DZ޽=u�xlWxs1Y�pG V���T���~o���z�8T���Ĳ	;�[�������ߜ�
Y���g���ۻ�����rK��n-mܑ��}�V,�]��9T���~�������+Q��O,�-�<�x����%}�p��R���֓�O,|v'�8��;�~s��XׇF��ˏz�xyW��������T  0#_Q�H4?��̩���:�3b��F���~����������ը�ޜ�WZ��`E01V��U��iEP����X�ٖv��k;�F[fV��n������4�q1�r��U݌�K�BEX
�Z�#��b�o�h�Ie��s05���R����}?LG�x��#�)�qp80O�W��{�������e��ǫ'��,��� �!��zvEk-"�Y-�U �5��>�;,�X-�gw�f,7����
A�@�j��Y3h����M�4ڨd����(f����"�v,    IDATNs�$ݾ��95V�h��ٮEl���UU1�On���N_����r�?�V P���H�bх =Ǖ��h�ZjhfHXF˪�D�����X�����֢�  �ZVZ\����%��%�l�pd4|�h���~�R��}��$ѽ��$Ѧ�-O,��Wx�j�C��O�
�!��B���-��BD���"a�J4(�v"+MV�f�4K�@� m!����r��z�\M�i�<>|z'�?���k`s*�V���bK 1I�( P�p ����#��xo���OW�� �_���o�֮/$ ��;P! ������Z���ok�Y�'����R �u}i6~n��X�r�����?>Y����Y��K����j�%�H��#��F����!��N�|p-����8]i�yj&�����;0|�����T���_8��ʽ��˰����w�g�3�s5@{�U�������H�_�H�]� `zY��ή�+sɋ�ˋ&�B�m�8_�i>���W`��>�>��/�����bd���+����"��/Z�6��a��_y��o�Z2���nme�#����L�Z�U���h�Eb(���ͧ�"|���������\H��ޮ����@�,c��o�̬�a�J��4��&�;ڣ��q��!V�fa�v"�M.�8P�D�D���x�W�@1�V"K�,�`�G)�f[B��u��?���(���JX�(�"4cQ�u��2�I��4�����om���/��ݯ^:Q^���[��w�^���������������RAa-��^h^�� b6ګ�!@�R�ĸ��%�+�b]+¾�,�9J$�P���B�P�0_ӊp�J!a-��q9�UU�Ֆ��6w�/So����h�Q��"��&w��5I_�'h�oh�J}~/�B\�#u��d�^�ؔ��Ԑ�d�&���o%�g����ъ�0^�Eߵ���4�����ҟ��4�z��X�Kk���йf����o,ڋ̹�'Z��? ,7y9u����B�Z.��\o������� 8��M����oD���o�Ҙ]��E6��V[줃���P�X<��Z�-�����YgֲS��NRs��[��! ��ϴ	+�"�]A��ue�*�~hc8�W�4�E2��o�?X/�d��r��mg6_��Zg�s"���JmF���vr���F��K���\�V��B�c�q�� *�5
(��Z����Ѳ�9�{�ٰ���Y�:�w��R7._M��"����x�N��+6��&|W���O��9$ " Jg/��A>!Z\32�����S��&�7�3�H���cK_t�Q��V��̝�h�+8�s��	���%� ���:� v�ܯ�*���R�;;�u�D��O��n�q[n�)��_�6h��D/w	��&���A)"�`�ú ^��a��|�ϰ#M�r�p]{�|4�q�A[iܖo@{5_�溅�<��v�����'c���n��#3U�A��Jw͎�%���4a9o�hh�͎ @�(��^�����.�֮AsJV���;@�-s�[ݝR!�f/��稆{N�� r�'^5�hPu��@��(�70(bؓw��:�	'�ף�n��lalS{EV�#*,�B��m�N�>#��ȝ���N�0�GRAT#=���J�� �K_A�4�n�g%DKVoB�����dGx8u`�'���F7߉�?е�[O��m�MC� C؃2���\y�hi���2�>ԧ��?�^�!� BBƿ��

�<ga�m�ԑ�ޔ՛�����V���Ij���i.'�3�Zܙ{s,�i�O�z+�P��U!�?��r̒� Z�Ɲ.���dbWe��� , b�`@Sl�g�Ĺk��X�~ޗC��K�d���xhw�"t��D ʦ�Y;P� �ؗ(�6IN9�"E`B3� ��\9� �9
9��6y�ϙbӸD�Xl�a5�MӜr�i���	ѴgG�ta�ghK�����9崣(d��L���=܀f����)���8S~gk��u�%�eL@Ă*��\�)���L"f��"&gS���Al�M�ټX�C�Y�F���YŤL��tq]TWD�N�P�E �d޶����HD֙���Ml��6����3л����n�M4��2����x��m��R�����JN$"�%o;T襱ǡ� ����3�?�N
4�, ;��d�ٙx�FOP���[e���r9m�R`�-��*����6��촭����zCnmy� �1*kr�Z"(��vu7���SJ)��#�)�K �5�!��gp�D>�rGlu�; An�!���0L/�p״VH������Y
� �� �0T��|�N�\���W��/b����Ō`�_A�-��lY����]�Ѝ��oҗay����=���/���8���g�gp�� ��զ���P�=�L�6>I�;_����
fz!_�/Ev?�a�,�$$@��@F���ͅ�h�nl�NErN[v�7]a$ڕ�@�rm�ng��3�����5s�-����4 �t�/֡�˺+Z���2������f�+�}���X8ԣ-7��3�j���#�����K��	;p��u3] ���Д���k�"� i&g��)�!�]�N�<y�С���v�}�ڵ�/~���I������D�T�V�533S�o��������j�ޞ={ ��͛_��yO��`zo��=Zz�@�m�2�/>y��槭�oD���p  73� T�oPE��Zң�jO��2�<�;�|;^^ێz�GW�Rf��ϛ��( ���c��&�@_�.�Ʊ�0_73Н�iF1� �kZk�d][M�v�!�u%?p��/�P(.]�444���0>>�ꫯ�������:�����@���v��/�˻/x���cǎ��O)u��)�jϬ��f�f3���GK��/������G���z�P���RC�!���>T�Џ߯�Y1CU��c�/��[K͑����\��<P����1ޡ��郅,�=\j����ȏF9�� ��G��}w��+sq��k@fz���I��"���TX3!���
����uxx��_^XX�կ~�n������?���o���O<��3�F����������}��g�y���/
Z둑�r��$���|����������G�������B�0::�q�R���w��������YZZZ]]-�J���D4??_�ׇ��}�yyypp�P(4�۷o���`�X,�J��_!�ݛ�6��>>�9P�n�f����ƿ?U��Di�����{ԩ��.5���B��ti��X����\}�� 0ңA�Q=ң�!6b9:D�,7�skx�^�jV����l7ڂ }e���i3����T
8\U�0_���P���@O��@ �d�yvV���m"PǓ)7a���	"z��7�����8>w�܁y��>�lݙ:r�����7��v�Tz饗 �Z�NMM�����zꩧv��]*����_{�B���hyy�Z������ǭV�?�A�V��ŋ�}����??<<����/~�ӧO9r��gff�^�z�����o~s���'�|���㸿��ҥK��w/d�����X��Wc-^o����
�c��&޽B��(�e��.�=\�@��[S3���GB������x�W-����m���]X�x���+�B���\�o����t��[�XK�@���q��_x�<X�@�BC���ƃ�
v8�#)� ���5������/�C�*hS;��ѣ׮][XX06' �߿jj*��O>��W^�T*�o߾}����j�������)�˓��'N�x��w������s___oo��/��k׮���0_�uf~��W��ǧ�����.\��駟����ڵ��ѣo��VgϞ���3����~V��qnn����;��αc�O�<��^�x��_|����@��3�7���C*�5+��BR)��$�Yօ ��Ӈ���o���H��GJƪLX~v����B���GK���Ԋ�<�7�G��K��y�7iV�4ޯ�)}x#:4����������% �;��i�෎�zK�� ̖�<9]�%�$ia����.�A��l�LV*��ׯ�ĉ ��#������V�A
�����>��w��я~411Q�׿����qLDa��Ap���]�v���+�� 0��h4Z�V��.�+++��ޡC�&&&���(�� ػwo�ټp�y�f������G�=}���ܜy�J�""���V+����6��nF|n�)d���ފ�����'��O, @�H�\]7�<�����I����׵sf��ppm!ik`��.�����GJ��V�A@�[��7�\���r�������m��T�uV1�i8\@�L1����3K,;���������|�ɭ[���}DܳgO�պ���T*��ݳg��˗�\�b����NNN���|��Gw_�K�K�.��������Ç����\�~��w�y��w���R��ѣDt�ܹ��%� ���XOO�y������� ��Br����X��╍��^�K|c!�s*��������L{�\m�n'���hb,�? �f)�T*`��	����������Ll~Y�d�J}e�-YCj��"pe>���;W�z�@p�t6 ���l��@l@O,�i�[���a7�<1`�=��O?}��'GFF����^�z��U (�J�Je߾}���w��>��}��������� $I��϶��v� ���A;vlaa�ԩS�����H������n�{zz>�����s��=��S���q���H�����C�^y�j�:77W��Ο?���C��a�h4��-��<��f�O���b3w>�u��'?��r=i��s���G�������#A������O�"��l�ߛ,�����N��d�c�_�o��[�����>U�����ZKZ�ȧ����z��N$ ��U}�z����{�X����t�����M9?���x��E�]���1K[�\e����>���������_^^��O~�I�={�̙3���罹���i���F=&I���Z��qhh�X,Cqnn������8�㸷�7�c�Z�8�}�63�shh(�8������v�P����0������?���࠹��,,,��DQd�ӯ��̃mN�FO��������S$ �Y�?~�61>y��l����N�����C�"�VCUUPX�x��,0X�@�ъ=%�-����/S��uN��� wjv�y!���GB�E��R�c-�%�-�P��.����̲.�_�@A;ٱ	���}����4I��0��D��{��"D؄ؘ��̉�X�y.\��j0))�ò��GGGϝ;�&�s�P�R�p�B���!1���)kL�����#����;GK���R Ͳ��Oo��	Wpw����}e��z+~��FsA_�:uOc�   (@`�Á�Խ� #���.� w"��om޼y����+Wr^����Mf����d�^��R�,���:k~Pw��gG{���["�u3�r-�@�g1�&��J!4� �C������GH^��es�&�X�����I=z@�/5�����y1���,v4���DAf %&$�c�"�b3��P d1����-ƯP��c������Z���r��%3��i�ȉIϴ���C[ЧI�N�6xn����a�������MI�t�w�c��'���+��p]�3�Qt��L�vc����H h�
#�I|�����V�+}��Zw��O�����;���,^��:o��㐵�'(v.��ulz��d{l��M�uKCR��u�]�r����_��~�4_���gv�%kN�-�?�oB�i�<�ґw�l O��=.��
�16@&
!H�q+�-�Q0�:�%�pBg�B9m*Ŷ�ٶ���@��S��2�������ŨV!B$@5�{�,���G@`lQaё�[�c("@�6C��� C�~[c���v�M ����PO��ށu3�g�g��j7*I;DP
�3���ˆ3����I�IX��"�$�v��Q����-�i�s���2]�w��c��H}�[X�[�w��%-���<�øY��εs�����X  �N$i1��� d#zȍ�*�����{�{)���
!�v�$�-Jgg�@ �v:�9�D�$L�<]����S ��>�.j���)���;�K�F�$_z�3��rN�5E�Q��<�]�R (��0��3s��>\��Ъ�������{X� ��%n�0��|Aa0�Ml(J��t�G�ŀM�A�r�����JE������z���:n�h���� �����g&�B�@�*���r�$����j�+q� hB�df%�:W�����Rl/wL{�P��$j �8ԫ}
�9��S�낸Q��ED@"3��(0�� �P��r$6�#�F��k���`� A!(��zy@I9��r�	�q�'Z-��q�L�8o(b��!��@0�M�5޴��N၀(D"D�y�:HV�1�Q������u��j5��DLz3� 
�X���A@8 W� v"��kBfRi��
"�"��A��du@UBU�3�%�[rz�XQq�T��t���Q�n}B>r���)p����	��E��g!@�N1��:�oPX�^��@=5�����-G$�k�v� L.#� ���Iv��+q� �L�&�Zkڱybz�:�Q ��E@va��KV�rC��`,�W����7 @��v�Պ 6�LE;ȄL��נs�vb�X�ӱ�m+���b�Pl�iӤ�L-� �q�}$X���� �>�0�Ü����)�A�A�u;�ۊ�L�"@$4����eh�LȎ��6�tYav6��(Fo���@l'�#��~a�@��E�$(��F0�h
 m�L<��{�F�k��IK����K��[�k���?��X��p��P���k#�в���n�R7e���|��%�� .���"~Y��L&���X�nw��]W1u⚘IǊ�@Ŏ�Bp襯q��ɮ�܎�ok7+@$O�K��0������c�� H�mpO�l�$��M ��wD �(N�0�HW5��fΌ[#�T6R����\����h-��-�����`ྜྷN}��u�c�%���f�b�]�݄,waz���j��N�a�hP/ @��L�s��Na��/��;m�`b������c��
ͽ���0�!���'`�"mm� 	��� ��鍒���$�pV깝�z�B�K!�H��m�""(@"�Z�@��P��V��G%]!��a��A���4����n���!��l��b	fVz`�G��b�
P�Q��YB`���[�DQ��@n9M���|VP"��46"t�w���G��6Vc�o����N<�O��M�K�=O�mI�+x��-{"��t��9&��]��Lu 0�K��kfe�k@%��-�! ;�h2 9e�̉���'�]�%�S�BΛ ���Zb:�;n�ؽ��)(�fO�<=��⟔M7Wsr��5�DȪ5LP���^�jIt*�F�\!�80#n�=B�R"��Ϭ"%WY@ ���,C
����Cڑ�kU��(A� �  �eu����+Y	j���&����t!pg�13z�o9<4?�����KVB�`  h���%v���hDY��\�����D��N�*@@`d��� "10�F���Y��{)��XQ��`F/�����\Ŀ�dXj��s�3�hs��Sz�ѩD#Y��6r�͜�K\��K��ЄN�ژ��|N��O�@7
�М2��h� !LP�6�r��lU[�g� � �n���6!��1�{	 �v�+V��d�]FCy�D�LY�;�e�+�I�,�ٍ����Ode�	&x� �@@@;e���F ��_��6T�ф�P�_��ne��e��R� 12  d�:�SP�����C�ā3���@��m��o~!Ȧ��Q��v��)΢J��gJ���b%^5��Lhg�|����(�櫻GC++R�1=V�A'�  IDAT��$@r�>��/7�	�L�q]���s)�F��{#V`�n/�3�E8���4r���FH&�l*alb"X��z%��+ʑ�S��� �fE�=�H��}���Ι� m�tofd]`�\[��|s2M30t櫰WmU��E "���Z�X��`��W� 9U��+��s��əqf4�=��sI$"(H��{�1)L�y~��{'��<�`���� �������2�Π�
��lM5��V���d�B�&����d.>���>� �� ���D�'��B�a�3Q��`�`����'HH�� ���	�Y�ʲ�gm2ˬ��AH�^���cɘ�� ��9��У$9���XO�^��M`LD�bLa�Y4�l��ȚG��mA@9�"V�� !�52ܦ�[��ޖ��)�!��b�5%o�cڋ�q�V8I�:�od��0g�Wx����Ҥ��Sga�16��e��ǒ,���[g�v���W�k�i�,p�+<F�_�=O:�ϛ��G��f��F�1*���&��ZȔ��Ͻ�ǵ��A�Ѱ4d�ɠ�a཯�n&�v�q/$59m�N���@�%�Yd�;������!dE$�
�p�U��A��u�K���w
ͷce B���.Z��c� ��Abf�����]'%������5���p%u\����je���	*4,��g�d�I�B�!*ΗN�$c�yC�hê���ֱ5D�8%^�Iʲ�`z~����0f����]�͈=b�a ��v�D2j�d�#��@���8�Fٌ9��`�:�����F�����l� D�Opu@Ϊq�P@ˎ�qJ�i���0���Z!�l
�;��S�6�ER{�$K�a��>�h�;���B�6�@���'�9� A�n�(���,��GeX3@+J=�xf _7/���6ܛ^�nxjZ�E ,��5;����dx�f-N+ �&�bz����� �@�7i��0��u [��"�w'�5�*-�;�1�!A4  r*_�(qm�]S@��z�؜�k�M^�{�.Ё���g�9�`ԵF�i	c.n���=杂!δGq�<�	m�x��(�XLE��۷�A�
oצS$��T��&R!��8gK�	2x�,k����=:!m=�̬z�w�bŦ[��рNu��WBK�8�'
�=��i��}�3�њ���II�-���n�f��l��3e�0V��h6.*�̘WF�5A��?���s�m'a���ˢd��F����
�mf�T#H؛.( $v�����W�쀀ʝW��id�  �BŴ��
��	�)��`�w,}x�4��L�@jB2�uMu0g�`b�XH}gI��T"fU:��'�`�I�K]����A�aVtaGo>X�&��EC�ԙ`���	���6h-;����t�-k��!���y7H�ya�.b,6t���"C���&f����p��3�H@���@�TSJ�z���-:8B��z�K��7'v���G���E���%c �@�|� �_/���u�H�f��3c਑�#>(�k�|q�)��7]7ѻX�FS�x@Ƶcg�zF&�N�I>�5	��d�Y뿂)�B�\ͼ^Q2��Ȯ&l��E>���Ѯ�A38Й
��=`�a��-��N��؛��b���W@��Z�>�cM�R��.`��D�
��+.F��*탊���f+�}\;I�Jtaq��?�6z�F���.?u�3�͖�̵��n��������吙��b�N3Gֽ���)�a�qn,���
��H6��-��`��X���S���k�&`��� ��
}Z&"0
g��8��A!��*��tI�!�����Q��c࣢B��ѫxt�(${pj@�����	n1L�?�SY .�@.�$�
c��:3��=�$���BTR�Jo�IGB��o�Qt���].��Xs��"�:�0�s�|�\R�aF6���������k"�� &J�?H�j�@4=$��|�ܚ�x�2e�HҬcm
h�S��!]�	)�&z��\\#�e�T��R5�g�����XVo�`��@���􈜋X"��S��a#��Ϡ:��ȯ���im�{����m%���Yݗ��dpq$v�:�h�}���fo X��
/�j2 ���)<��E|�'�dr@d]��3D-�e�ѡ�EA4�wn>)��,Ȑ�p����C�?��+R|U�(��[0u+���Ƃ��В
A�@.*��jƤ7���c���W�n`� ���H�HS�!Xh��FIr�(R��^�Iv��/�2)�V�X!�k���L�׹�)V����uc1��5eI-{r�")�,>��GŇԭ@p��$iZo8��"��!����S̚�5��UL��x���o������[�fkռ]�`|
�y�؄��%�y�˥S���>+ʉc[����h���{�eR��u��r�th�����un�����m+��Sy\���Ohԉx��-SY���"�!p^2c�3Y�) �ۀ��ʺ\N�m�@���^��i3��?޳󈭇����a�G�A���aZ���צA�:�l��[y��* 
3x��{�6���E�&�%��.!��2{`�]L��7�ϭ�5N��{��\����'ٺ&��
emn��b�sb�.2�����5���9�ƺÌ��:6.��'u
	*��H��Ko#+�]֖ɡȊ޵�F�I�(IM��Ku5+���-RC�>$��=�<8��'��8HU�!4w�=p���g�#�I�2:?��{k$ ;��j�l��-9@��ه_D��:J�/|���P�@(�$RA���4�-��kX	=禵x�2������$ͫb    IEND�B`�