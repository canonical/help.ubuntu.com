�PNG

   IHDR      �   �EP   �zTXtRaw profile type exif  x�mP��0��q�8N�Jݠ�TIۓ|<}Ɣ��|���"^�ޤ5P��ԡNǘ���'jzx͗��@ ��aon1�q!-���P�Ga��C�	�Cd�x����U/`�4����$��b���~c^u{���P�	�2� d�
uHYk���$��{J�7�oZ4�]�_  �iCCPICC profile  x�}�=H�@�_S�"�q�P����U(B�P+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�F�iV�,�鶙N&�lnU�"�D0Qf�1'I)���{�z�Y���}j�b@@$�e�ioOo��}�(+�*�9�I$~�����ό���<q�X,v����dj�S�1U�)_�z�r��Uj�uO��p^_Y�:�a$��%H���2*��U'�B��>�!�/�K!W��B������w�Var�K
'����B�@��8�ǎ�<������W��'���;����붦��;���!��+i
��~Fߔ"�@��[k�@��J� ��h���}����ۿgZ�� ��r�(˞�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:11a37ca7-9760-4dc1-8aa5-0c1749ca975b"
   xmpMM:InstanceID="xmp.iid:d49d3b2e-99ea-40ca-a0f9-633f30b2af90"
   xmpMM:OriginalDocumentID="xmp.did:e738023a-9ea9-4cef-8c02-03954f0d3515"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679601694177475"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T21:01:34+01:00"
   xmp:ModifyDate="2023:03:23T21:01:34+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:cbce2f3a-99ad-4846-afe7-5ef4d5481c78"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T21:01:34+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>�!�   	pHYs  �  ��+   tIME�
*==   tEXtComment Created with GIMPW�    IDATx��y�Uŵ6�V�>�9=w�̓������(ΈS�jԫ&*11z��3�Oo�����ԛ|�Fo4�c4ƨ�C�AQAE�f�n����8}�a�]��?j��t�>=�m�OԜ>î���5Ԫ� 8p���88�t��A���������^���B�UaF<O$�tZJ���`Gqqqeee ���i�����l����N�������C��|���ԝ�|�@ �N��p$�������aÆq�����/���@   �X����1��.�`�֭������N���ٓ�c�3�	�nwUUUv@ii�]w��v� ��.^���
�~UU�̙3/^��9�(���,++�D"?��~��_꺞�f�Dw�z�������Fe�1g\ bEE�bN�����x
���!C��iӦ��9r�I'����`0��o�駟>��~��i�<���~���c��Ò���g��Z�������.�4����떖�/n��3f�?����N�2%�H�����<f��g�}�嗿��뵵���_|���d�y��iZ0t�`p�^��ǯ555]q��}��?�񏫯��G�����'�X�x�\.�z�N���ÈF������������/���_x�D"���X�nݢE�&L�p�g�i7
96��A�c�.����?��s�1����Ƚ�bŊu��uI�3fv�e˖-\���tIIIw��|�1cƼ�����G}Tɱ͛7��9f̘�+W���9tfXw���M�8q���;w��f�ʈ***=z��m�6n���5�䭮�7�+������ڵk��{�
���9�R
!4��	��K/m޼�駟��O~�w����s����������p����?�|�ԩ��p��g�ر��<O:���2�L}}����z���4i�|߾}�mE���hv0X�W(�iV���+����;C��̙3����]� ��o���[���Y����;/�T*�nݺ�˗2������v���s��Y�xqkk�ȑ#��x����ϟ������"�p�\&L��w��L&_x�Â6:#���:����a�d���w��q�7t�P��\�&M����q�ƍ1�;�����SO=u�}��7~�a =zt6�=x�`)�x��!C��}����ͫ����g�N&����/b�Xw?B�>u�`P����piii�Zb�"���.��{��}��'g͚�{������U��<��D"�-ڹs�y�,X���{･K������U<�i�N���A�������#��f͚;w.��0��˗oڴ	 �:��O?���ҥK�n�:!���ݻ�!����yuuuEE�W+ҷ�����h4��DΠ:T�b<7M��vk���:�����ߟH$q�8��`����B���"��3�\���H$T�Ǒ���^����,�T�����~��~��@H @ �H"  �Dd6U���R"I 	��P  ��+"@� �@`_��>" !#�B@@ @�8Z7��[�$u����>R�"@@�.�T́uod�t���'�H]�PJ`����@]@""H @�R��D	�d�!H�$ 1"��������$I�d��՚����'�`���5#�H@���	�@! ������ P=����	`�!  ����\!D5%�^���W ���K��]�5��H�|�|�=7<@��S�@ �/Y�A������$��n@�˒	`�$�f��A�^�jBIi��V+Z�W�@H֛	swH�j�#�}�L�؁OII� H���	P"���)#u! F��^D 5�C�1�y�nB�,���>!1�ĀО�j% �dVǒzN F@�TϢ�Xk�H &�%J��H@�Pk� �]�t���5�A�}C����.mw6ؗ��O��Cf�Z���C�% S1 R\D "i�TOl�"j� "$��zE}`qL�k�E0Ǩ��g��V��$�t�,IiS�^r;H�PJAR�a��C�9m��>��˭�Q�}$��T�( ���=	@� ���ڜ��[�DĬn�ؑCsDH�T� �ધPMU��N]�H� �)Q$�J��Z�	�^' � D@֬T�c ��� Jbjݒ���$�M��$$&� ��k$ `j��5�%�$ Jk9�@�I �s�NS���E��IB@�����֘X�'��G�-�mY���/Z�:v�����"[�Y�/�PZJ���BHI,��FT5�vG�P�ڹy�Z�'AN��2ז �S;(���H*Q�1�����"  �d����5����~(�^)�����Lv�K�T���,t�K���Y�~B��Cb[,��1 P�U�H9�M�(�]k�E j]�$�r(@�T�2$)A ���wK}Q�
 � R=�R�$J��ĉk��BB)�h���1jh"I ֱ��5��BɈ���aNP3L-�R�N f�ˊ�?QZODL�gѦ������JK���	���`}_�����P�1�i��)1��ڔB���� �si��HJB��K�Ԋܢ���A
uyKw��\�i}6)r�~5�}!�RvTS�$��|ˉ�̭\և�1O:�P-3����E%���^[�6�����H!@��7D���)��Щ_l���/��T@B`���җ,#G�J�D�d�� B"	� 2�E��Ą��dY�L A�:k����ί:��Φ�!�#[�����4K�8��#����:�8�(��;��Nd'c���=�m���>t�c:n1�>��N�JtؓS�T���6g�vzJ�.;��ut��uѝ��TZ���n.}��׭���>�_�0��R$	R�`��`&�Q�*Y���Jd[2�l���DF �i����e
K�oP2��4}"RJ	BH]PpM6eZ
I��8�G^��=d��i�B���1D��<�`�̤�i*_*G
��1u��:|��)͐J F��"(	��Y�(I�dJiJ&��lwV6�"*��0��W�9���cEŬ��:�ǡ=,�P�7�|C"e��~p[<�F �s ��CX=��$@�)	��&�SlgF6�zZ����R*�����R+.�­����W��B���l�v��-w�e�� id�pW����C-_�f��j���f�� !��� �&��3K���a�Ս$%���4�&Œ�#!�f��|���/�G�њP2��-�O	5�7O-ϓ�#1R���ъ��$Id�d�t0�b���v���kL3���6����:��)#�ٟ!�{�d����R7�-�6'��T|�5F)��*��`@Z;����f+�����۴FD"�@`
0�4tٞ���lS���8��q�%$k?�yC1�o��Z�|*\�ڄ'�$�0e6�jRF��.��|TTb0vЖ
d��H�� %��" `@( %�d�2�­	}��0t�k9F�����Q�X@X��v��@�\# @IR���0�9%�v9p��cDFe5g<��v�1Fh�%R��rlHi��J�v�L9���A!�AQ\�bgUD:2R��r�增	�$�RY�7kD�fz����{[ёG�d��l��Q��\ζ\D�Ѱ��-)Ͳ
w4bJl��%�4ȅ}H�ڐR
cj�r��4��T
���aH��l��Q�J+<��P��Q!��9s4�""M��%,�j"��@�fմ��I��f�5gE{��@D���9�.E�z�s�9B����X����9�y�F6��i�X���jK�����v`"@�>�cD!I���+��s��tQ����a����e[�*��8�4�s�3M�0�A�qMZ,j0��iX�&��$@b�l/|��{<��g|g�tW�f0��ਲ�����A�h.n����:Vm�`H}]��@��au��,""����/�X��B�4�Aؖ�c ���sM�
_+�e[D��!�ϭ �S�H)Ȕ�5Y�@m��w����\�X��ਢ�+���*p�˶����R!�$%H)`.���!��R�j�;�<��l���cl@�B2�˶r,��@GB-��2� I"����B�/���Q�Fy<)�={��#��4�<V_�m@IIɨQ�ZZZ����wV��U�p�ͫ�2����F��L&������$RJ�W�Y����ї � )H
#i�/�Q��H��{��W���W^y��_��xv�ؑ�d�Y���y�b�UVVf2�뮻�G?�Qyy��U�***t]��"ǣ�e�����s>eʔK.�dҤI�H$OIE�<��Ƕ< <�裁@����s��/�`�Hģ��!2+'0�ҖJB�dA�N�N�<��o?~�������t��O<�����Yg�U__��+�|��GG>�r�v��-MӮ�⊫��*��=�s~�Yg=��3�@`��Ջ-�~a��m��)�gϾ뮻��s~�<��---����8�qrΧO��p��W_}���4�~�핕��>�l����3D�i*���tR����V~��
!Xww�wTUU�\�rѢE���s��B��׿^�t)c��;�,**���|�r��;#G�x≈�k׮d29y��ѣG��>���tpTѣEt�7�޽���~�G|>ߥ�^����'M�t�}�E"���Z�Ά&N�x�����>߼�.Wu�0�$Zu���D�'���	&<����ڕW^��o}���J)�}��g�}��SN����Ds����R;kkk�~���������k�ԩ��!�HEg�)6X�/:t͚5---����H�������ѥ�^*�|ꩧ�R����?��sw�u׬Y�V�Zշ�WL�P���sQ����V���=M�t]2d�u�]��{�]���<�̂�N���f�[�&�~��̟??�;��k�֭khh������~�DN9唇z(:�+A0��3c���;q���.���K/-++>|��	�v�<��3�\�l�r����+�ׯ�R�]�v��ݳg������Mbvu���0%�p��"��]RR�iӦx<�aÆ@ �8��3�<3
E��p8��T�x<�L����~��>�o�up46~��x����}��g�}�zsذa���m��6�s0������-�
���ܻg�\v_��ʄ(U����C�#���~�m�]~��?�����S__߷;���O��-[��3f(��s~��'WVV�۷��G�D"δ<�3gJKK�vc�&M꛺������N8�0sk�Сuuu�}�C��#��/�v������}ѢE�D�{�6l�����v�)��]��?ܰa"Ο?��;�?����z���{<��;w���{]z�,��`~�<�����f͚1cFgo٥�^Z]]�bŊ�y+�/�hz`�I��D5G�\Z�N��g�!ğ����^{M��dN<��3�8�������� O[~����
 |>�7���.��1��͕����a�`�RʁU˳s������G�����W�Z����|�s�=wҤI�=�ܞ={���Zb�niva1bVj*�`B�.ॗ^����;�#)����ꫯviI)�{ E�.�J�Ro��F4mjj�袋&O�|���?���UUU7n�N?<J�d�!Dw�L&�J���#U��,O[�p��g�iii�;w����/~��_�^�:��[��QE�:t�o��Hu��0D&�jۍ��:pλ�w�\%%%��ȏt]�D"�l�ȫ麞g�������1��sϽ���}��_|Q��]g�o���C��|�����H'�a�ž��٥	�c[��ZTT��z�(�J�b�<��֡�z�o� 1`	�g��$�0�Ncm����H"��; _J��f�mǲ-G.��ǰ�u(��9H��D0�E0dȀ$uk����!���L���:ǲ-Gi�Ǧ��ft�|��  0�TxX��BU`�cٖ��"��Z)��u����i�W�*�ۅ~�$����@�t����e[����?ke�hs,�:�e  ��	��*�{��o� ��9t,�rpTaF�;%�z��˶:؅*a6j@*�Cm����7��ʠT){z��ǲ-G�cj��s�cٖ]�T� M%J�=}
�P�^�<�Oߣ�����˶m��B%J��"V���}^%�Y[h�'R\C���j��j����T�3r��V�LR{����ar,�rpT}���Nȝu��VC��q<Vm)k4 $��MP��oª�X]>ရ�Ǭ-G9���C9��xLڲ0 �$�|�b��Z���*�����O��*� %Z�{�7:'8�d �8!�*$�(p�`@����B$D�p���2d������:p���כZ  ���F���8s�`@TDBM�9+A�}
�u����̦����@�-~9p�O��8 �uD" 8�8�/��Nˁ@�-��P�Zq��A�8���D������L��Á��Z` V�D�r�ˌ ��kF���Ǘ��}��GN���`08iҤ��J����kjj���_a������^H%����0�ǳ`���_}�ر>�`,s�#�;��n���O.))a��b��[�>���6mr��}U�0R�ۘF��	��XZZz��wWWW������?��b���/��Ώ�ӧ���?1bD���s�N�>��\�r��E_A���H"�*�h���馛.��"��:��<���}�G�5��i.�̮�J㭷ު�;��ꊤ!���AE��|����>o޼P(�r���7���o��d
8��_9 �����㧝trw�N�0ᬳ�z����%���0�~$̱|�����Z���K.��s��3�8c�����n�mar�����'��(N85����\S�Nݾ}����K!X$�v���-D@�\�Vr��{	���%7n\��Y$y�����Qd�d_�Q�z(Y[*�A�fu߳#���F�)�!C�}��J�ӟ|��)���K,���>���X�ƧX�䯧��n�y���uM]�0���������R$X"�菧Cm*k�P�U���H$=�PUU���>k�, �����3��b����y�h����Oꋚ���q��u�iSS��ի[ZZ���Ucg�>�G] �H2Ml�PSo��D"�����g��; ֬Ys�7�?���?O�RN�w�l6���~ꩧ��}�hѢ<��N0tl���2�$$�R
I�`��l�N�Ŷo�>jԨ�^z)�^u�U�����lw�������>y�d�ߟK!�����?��꫆a8]��#X�"#�fί	$I�"�au�bS��V��ٳg�3��_t:�G���]x�&Lp�\{��Y�dIcc��-_Ep�۱�d�9ë�<� %H)t��fX]d ���ז`;�
�6�$!:���� �P�O ��]:a�d�J�#YY�PEJ9.8 z!!�;�Y�{G�9p�O�:u��@��v��}~9p�_���@��R�� �`d���	���N�6�/��yBf�UAˇ(�9p�Of�BP�D0Wx�`�	f�1 �8�� ÐԎ#�:����A?uD[�!iJ�媭�3m o)��c�4,��Jм_��!sp�T
C����>�y�ѶC�����
��]��aX>�&��\����&�&�Q��S�Nj�J���~눖��uT2R���H0>�����c�i_�Q�>�y�K��Q��'&^b&���?N�Zj���l�)a#���9�|p�à�0+NX@�Vj�T�]Fm5����O� �H�$i
����%0V���z79���b�u!g���'�8�=l:s��p-���3b�N���G������Û^����qXux�)��L���6@@@Db|���<�$%	��g{K0��'^�O��8��G�u�,�z1�u��&'26�m��X<�k�>��e�
��ɬx,Ej!�%�\�6@����^Z�V��S�����\gd��c�,�u;���]#��o o��{Ƴ�����18���!"  Cd�A�D����46n=���    IDAT��M�|�x��2�;ⴢ��Cw�"1����A��v�r?���ڱJ�H&��q��&\��(�3�t��9=�� ;��)qz쨰�b2sQ��
"*�Pc@��*� �q""g'\��a�%0�?8�J��AE��,�t�Q����ez�Be�!i$A���B�U<�U���׎�r]0��� 6�חoO;CV8��ў3S���vCq���z��$C���>]:��b�j6|�8���R^D@M�,b����m0d8�t��z����o�)�ژ�L���b_��-1�����gN�yq}��z�MΠ*��ERrX	OԞ�cA�� �Zb�̽���95�����v��G߸sR;�at��`��­��gi�Z]�-�w����<�F�MhO�d� `T�M�h��e*Ƶ�TG}��n�
�}���G�[_��Z��S`HĈX�io<EXz|!�)G���]�x�/?���e�}]��o�|�겇/+�4�}�wF�rD(b�����K.����/+���>z29����s~ѱI�H�﹠��!���k�jW��n�ۃ品�l׭�����<%�su��}?y}�C����ue��_����,�?�g3[�x�Ɂ��݅���2�ڙ����I#ܿ��"��;��-Œ�
�#���0"R	p� ��.�.�@u!�l����& �3rgK�i4��)u߫��'"������ڨ��,��bxУ���үmLni���?+�1�w�@X�gE^� @��B^�V�"/c%~�`i���L�l�P�c�~�/ ��2�;]�����n>�,����s�F�k�����U:�[���N	|��?C�e�����o�Y��^�����h��g�����|�]cP`�A���8�QE^��t�ic=�W!�ee�t�P�W�&V���Q�ݚ�܃�����=#α��^Hf+u6j�{	$�����¶\>ؙY_�]u��ǗD��ڵI�HJ�.CЁ�8 ���A��lmm6����^�{��ŻѦ���Y��O�K��__�U#z�Dבּ�������"����7��T�z��oo��k3G��d�~�}w�y��msCǐ?oЕ�x��Py�gMzzEl{��­��_=�V��6��CE�����c^ѽ�ϲ��f�;�
������=W苤��3C�*4��͝��8��!�1��r�2�X�j&2���J�/�-���0C���?�{$m����xƐ�^�X�]����A����g���ӂ�~���<Vs�[��{Aqe�gMz~M��}ًO��كJ~�^L5��%%#J����ǖD���,bpx������T�PvX�ND������×���u��'�)���������G�j=*�>7���o|�\W��Ż�_�Y�����f�lI���xsL�ܟ�7菿m���f��t���miПZwkx�8O��7�
~�l�lqdW�	 ^��)~)�%�HJ\4���0�+�O���s�|ze��񶹡� �g�|�~T������Y�<��wc���q]���	e_��c<]Zrͩ�+C�ޕׅW�d<�$��҅�}kk����?����.�w�-sB[�ǗD9�o��5���`ڠ��=���������e�I����m��Zw��q��u��C]�|Q��Bw�-�K�UiG�F:gLZ���I��������ʹN�ʴ���i�ztd��&�/2�11�T�����E>Vd�ʵ�.���l;���eN,4FĖ}��̸*��;�a$��f�=ٽ͊ ����ek�{� �w���ڄ!���.�XK\r���6�"8��`�!	G�@"�x������XZ�����{��t��4�V�'q�~v��ck\$�RI˶�^�y]��.��>�~wf�W���)����lmԗlI�,�<F���i� �0is��am6cR��|.�,O" i�H%�AY�ii��W���G�;sCߘ����3�O�9���yٕ���1����][ ���Y����%gïq����hJ
AP�g�E#��� ����tIڠXF�i3�[�d�̀�dW����Ei�~�*ޞ�^"IF�ۏ�4�{��?����B����L����ڙA��\�Hd�k���2��oG�|n�u�)�:�2�����⎎"	ʔM��Ѱ2��)�ZRdY�1��eZ$-AjY��N�� =�h$z�/��0��F�@�P�B�9�e��=�~u}Ō�n��[�V�����9���U�Ui���w���Jh�ݤ��8m�'��� ��Vs[�������rm��z�y���Qe���'t�>o�g��Ͽ��|�%��у�X�E�ڙ���z��j�Z��.��Y���-��%%є�hw��/2GC��-�8��ǗD#��E�4D���� �=̭�?}���'�WGW�ޕ9�J��$�����]l�h�\\Rd�A�hU "��I��������K����S:�ms��s�~��$����+wf�6�L�e���Ԛ]��g�.>�_dO.�E���-�o�<~��"��ؔ<��^�8����EŋVſ'���z1���5�!"J�V�oa�I�(%�04��/�)�\��J�c]tL�����{��xG���D�6m��4�$LJ��'�5���d")����;��<�4�� ��Q�Pd-���}�$X�-�֥����"�e䯗�j[ͬA�,��J"xa]bW��ql��>
���d__�eM��l��r����T<; ���2��s�ci�����H���̘�{��Ld)�K{2���dne=o�ϔ��x}�����OS�K8 l�Ou���F �Z�2�����=����>��"����Բ�l6A�(��Y�g ~�A|��l��v��;�X�Y�`BV�XcTlާ����_��0DK��O���2��ú��s��K�w�C$���k�=@�H
�0�)��?�
2vµ|ҵݝ�x��CF�i  $��r�ǻ� �޽C�הt��Zw6���*�1W��줡�+�~�&~ *z4��暃�����0dc/�'xA�����z?�ꋌ)�h�� �f,�N!��4���p!1�!�\���
�MO���񗀷���>�+�%u�k���^�
q�'֥��5��ƶ�=��eݏ+Q�J(0񙕱Q���	������_^�XT[� 5 fm�!I�Da�F�Ȧ�٘��<[�Yv�_>I:��;�:\�mؐo�M�5�.d��}H=L�D�lX�kG""1�'$�)�o�BL����;p��~=��yC$[{�ڿS��鮣6���E�z�.K�1�:�D�
�~�����ݗz�f���ԯ���BzRl�3�:]vT�ÖO���� � �1 $�v��.m�r��b����}Ua����}���tA��a����cN��0ȦO̍�#�;ba�#&Q�$�V��ڿ$w�+��z���B�ny��Eԛq���b�96��j�D~���j���:�&�ƀ�l���t��;�Jk��[�x,h^gl�:�Ҍ�K�\���6���I��]
��'~�'�	�qгF�8@{�u�A��c)� ȧ�] HD�$�D2��y� �*�7B��E�-�]�:�:m�oL�Z��bv�G}I��F!�.�6B� j��9��z݃�fڷR��I�_�/Y�sGr ��P#+lJ���_���A��ٰC�r*�%j��aR3�z\a��.��"�/۴��l�D�7����_&�G�O²��D'uv>L�l���)n=އ��Gh��r,h�Kۆ���B�Q�F����RD���@O���H�.vt� UJ�����L�z�w��AwP#��"1� ��/�<�\.�\�_�OE�q0�*����r��A���󄚥"Z���r��:"S~bf&iJ�D -�с}�;�&�lB��|�b?+\:p� ���V�l��.M] ��+��ٲ9�1�����aB)��B�bÊ�X6}N���F��G)VOaU����5���ν�Tnz$"�]7̀�5MS�rƭ7�0h��hf����K��)a#��sЩ�����)0�bJ�Q�r�����@�T��HJ!L	}ι��r������4M�4�"�ǲ�ٔo��㜐�>���ǜ�CN��+�oB���J��t" Y9��*�\.��i�68 4s�\�hF�8������p�SEv �W�'^�JƋ�Q��O�	R����fGKa�إ�32M��nw/�5�O�W�]ɳ���ɷchX�	�FH@� �doC�4M�4�L��C��q��8�Osj48�VN���cj�.D�ކ(�H�Lud�Q����j4;=vTXV>����W���C@D��ܠ$ I {����On�z?�_��GLc�.�U��\r f99��Wa�9>ã>��)�b�c�CO��:�˵�=C��.hg��a���J�{%L`>�5�;�D�Iճ���Q`z_���s�̙3gΰaÒ�����W�\�{��#Ss�9��v���L����+--���L��XQQ ���_��j��-��rZ����$�M��|LJ��n^4���V�7�^#lh1���P��5UE��A6�D�m5'V�v���l.��?�\�ê9ש�!E �cb�0W,CBB�w4�_�$ވ����zsҙ�� I "S�bo��A������㏿��{�=�܆������:}��.�(�޽��/?��S,�5k�%�\RTT�q��#/x�5�,\���7�<6���z��SN9e���_��v�yٸX�m�`��[g��*�3�����^h��bL�Y0տi�>�f�#��^6-�~wVpS�=vUyu��6;o��3�u��#���0�Yq���{/(~eCG�&�����HG���痜:ڽbg�Ǘ�y�8��u�$��{��8�`g���O
�0Ř;��BD��Z��
BG��BV��쪬�����_RR��C�۷��������ZWWw����z����|��a���w�}�������?��_�d2�`��r	!�ɤa���^����T*��d4M�B�˥�z"�  ����;.�+ b2��u=�H. �d2~��s�~KD��`0���].W��/�c�u��S�����g}v�cH���lCD��KKo�|��a�.����}�$ ̝�U�m����]�=mF4-|���� ���!�C�TЃ.������")���h>�"���Q!A,۞V���B��A"K� 7ǀ!�%�Ĳ㩭���O4�		�h O�̝;wܸq=���͛�nwyy9"�����W�z��.����۷+&����B�c���.�N�B����'%%%����曯����3s�n�喙3g�6<�쳥��?���F������C�����oܸq�dr���+V����N;�4����'�<��ӷ�r�ԩS���qժU���7C�P"�x���w��u�E]{�����5k�|�Cۍ*�c�拦�r��:�������������p���+ĳt�4ߒ�i8��=i��j׭sB%~K��|�do�{g�&uq��6sG� ev����I�f's!`�����!���<;8�L�j�nM���!��Y��#ܭqQ�?{;��ٸ���ic=?ڝ}jy��08�`��,���%�e�p	�� �3gΦM�jkk�} Çg����w�y�[��Vii�a;��sO=�����/�����,�>��s�lv޼y�_~��ﾫ�f�ҥKW�XQQQq���Y���������)��ٳg�̙��_֮]{���ѣGϟ?�w�������_y�e�=���uuu�L������|���=��󛛛��7�X�b��[q�F��n�޶4�~V�?\�T�W��9��-.�b |n�yvpw�����g�n<=��Z���zy��՘5��,��_����p{J�3�I��}xx^��I/}��N�~fp��̴�3�{�K��j�*Z;��u��oV�C^v��K����%�
j~u"� L�DD�.6lŊ�d n��eA����n�;���y<���z�W^~��ɓ'?���\p�[o�u�YgUWW����v�8��wܼy�٬���  ������bW\qEyy�ڵk?�����;�s�y���].Wyy�W\�J������xSS����q�ԩW^y%缼�������ZӴ���o߾����+��ʳ��?�-1sm���3� ��;�K��������e�4�|��uNH����b��4 ��	z�u3�o�4DL"H��R�E�4�3�x&V�4�!�=8�B�����AϚt�) Q���U3i�j[L����
R��$#R
b��X���d2\. lذ!�}��ǈ8f̘iӦe��.k�I)��ۧ��	&̝;����z饗r���]y啟~��c�=��f��1 0M��'�|�G����ϟ�N��������?���MMM����/�0
����-[�ͦiZii�r�nI�{����[r�w8)#]Ն^�+���RU���A���b�9+��]�L��������#�4 �\K����ʴ�O�-۞����$ ��N�!�5�daK\&=�a�Go��Fx���+��I.E6��0  �6�
��@Dy�ď>�h�ܹÆ۳gϒ%K�-[&�������ӦM۱cG4=�'���=ztuuu*�Z�r�i���k����r)?ukkk(:��s���^8iҤ�*qVWW���?lnn3f��իkjjV�^}�m����pΟx��7����s�̹�{Ə�}�����6|��ߞ7oިQ���gsAD�����<u��@��f��)�n<=��L][���}���&v�6�Ċ�kf�<�[�Ϯ�Y����ǉ�h�缢�.�li0�9��١gV�3&@}؜?�w�p�!���DV�&		����y�r"P��w6�f�W������+�F3"R�Z!"���/   IRJ��'L�Mp&���x<>�����5k��:�$�8���<���_���>�<o��dCC���kjj�|�ͺ��x<�{��u��}�駵��������MMMk֬ikk���Y�v�]����՟�t:��ܹ3�b�D"�~����?oݺ���1�o۶M	�ݻw�ݻWJ���������U�V}��555MMM�v�z�����:K�/�]ݞ^A��	X2���&� O�V�l���ݚ��q���+*���oi�5~�K���8�)�H%�v���퀱�]4F��6�6��%A֠�VS�}�����z}_XD��@Tl;`4�D[BևMS ��HRֶ��벭	�q���}W������d�%DCD��t-ߑ��n~�`4EE,-k��^���'H���"w<�F�V���#"SJCȬ�m�x�"ӳ��r)�;��{&Mz��';O����9�^�d2࠰M���
٘�����s����'��=;T�Aiwum��Vŷ5��=���p�4�i�<?�k{[b�N�Kn�f "J3t���G���8 ���Qh] =�~!D�H9!�ҥK�.]z��K�,q8�+䉓 j�Jɦ<����ڜ�X�O�*�I�����zZ,ۻ�!~�9�����>9�E$�WR��1�h�BD͊J$Ĉ��� �^�|�Y��-���3��O6��U=�h��n�o7�36��S�bK�t :o��eÇy�,�\����P;a`zz��4M'��˱�:9:d�bvF���ACPCD �AzҔuK(��0�1=�HS.	H"X.����9#��c��X�B��m��I��e����Z�Z>�{�� �উv5f  �� c�dJ
W�L��u��u���N��u��g ��hXr	y`����� G�lF�C�Ș��U� " '�Hr�~���Y��]�z7׋��;rl ����܋�<��H�����||��� @�r�
OЧ�S�gl���0�O!�D����)�+�[�dD�Z�8@;_[��L��1�E��3d��q��!0B���$ Do̔���u��3J}�����d#�y#$����W��h�u&��~��yI���W5�9��/w!r��	4 $T%��#D�A��s�R�0  �IDAT�cj~�#LN���&��Q����_&�c��&a�D�U��I���R�lb��)��AO��F3"2t��] �x���FV�X$B@d�L$N�*WY�4�u������Z0IPd7Խ�����Z"�&Cd2 $ ��K��90dH����5G�w�'�%Mo"�"@K9T������*���#�!j9&�ܢ�3�t�ݱK�<�6�a�$��+#=0$b��,!!"Gƀr.�u��cG9p�%4�%��lJS��\������K*)pDƘ�э�EF���{�"�c�.͕J�a "p���
�@Dd���}:Ye� ����!0̆x|�Gs��٥�_�KJ��!rT�_���Y9n4��%�HD�H�!�HJ��
F�'T�˄�t��]��2	{�[J�"�Z���2�-�Ӏqp1t#�d�Xl��*G���?�W�{��@��-G`m�ʈ�������_+a=#$`�p#E=�-F��)�oj�v�|ݨ�'�=��I'5"�0䄜'D �9m� ��,zH�jA���B� 4I�HJEFi�8 x�N���	��;����5SW
n��R�T�`K)�_�w���ل�׃I���3M�D !	 ]�t?�ĵ`���)���9p�ՕZ�ٴ+r�m�H�K�Dij;��PC�#D��� ���T1)�C(�# "�12%�@)%b�C�|1�ň�%�� )�o��t�Ŏ�Hh��J��d�:�j�GD+��-���`h��h��%����_d'�%  �T�>d�P��L"����@H�2�)bZ���R��A� 3�	@ٷT��I�v���A�:F7�	9�l���4������� 3u����r]�s!,)e3�#2�ߥ\�)_�5��C T�����&S��*� "r@`@ q	��  �.2�2ňDh���l%2suk��� I�jB{�@IT	v�+�j#�l#�RiUxY!)�I�AeP�@�5(��(�Qϗ*�֭[v�B�z4䚚�1�DdU'YF��D"@��ˀb8${S_�xdU?��=H��.N�v���D���vF0uiĝ3�UfT�e	���&�m�2Ԁ ����2'�NH�� #��Xm�@"T�j=R������@�:�+swA ��)��#�^Z��$�DDH�sС5�6a7�&��eV����V��H��Y~�\ 0�v��ܼS	80W�!7�T���F��Fu;���������8! �I ԀJ�<J�����ζ"H�'AP�d8�+ǲ�K" TB x�B2�����h/"�  ��BB%h�L`�LT��!i}�^N��C �4`�[�<T?��Ȭ���H�F��Z#��u4�v,1+a�JOО�+H@ &�,G� �㠵� �T�=�]�^"�\�#� ҪlO5�C��H�a��.c�G(U�82�׀H���z�N�J��b(�m��G�DiQ��!Jf�)���$ n�a(Y�<�I�]n���ZR��**P-#��#��$; �v�3D;
�Ľ�f�� �h�&�ZQ a��	�m�YROZ�(#`��#�z�$I `V�0#d�Ԙ(���۫��=	T�M{A%��"J�� !S�yH���I���P��Ek�I����X����[m���ՕmK�� �z����vd@+=�w9Y,E�$�ʧ��Bڨ~��l/dǧ�ǉ��(��^�u����qsC�S�n�GH�cC$�sk��\ �i|ͦ� �=KǄj�}S��Ft��s�>�Q� [T�[��X�F��6X�d�[@i��@����m\ ���=��C�w�h�����l�-�qΑ�̳���V�J|n,u������6��d�v%��;���M���/�{%���8�R�a���P�%�`��� D��B��	sA� ���U�̔��i��M���b��.i[#�9�[J$��p1�1�����׬f�[��i*h�yr�MIsnU��!Ī�{�3��JhO!���K8�i�Ҡ�\O����,u�x��&�4U���%�{Cĕ:
�d�9�8"NMJ�9����W(>;x;��M��i�nH��Ɣf�'��w��I��Ubh8��C�����;��0�[C)����+���.�ϔ�c�Õ�ڭ+U ���1�#@�2t���*O��=8;��mD7	��I�xTu�B5&��4E�Ć��@>CG9��*���)��Te�nM��A�9 ����&�e7F�R�\�OZ l7�M�!O������9�T��H���㧠�:�%�b�ND�A��H�K2��j�#�Ul�T��:��3Z�'Iݐ�H8��q�הU�B�t��
�1�Yd�/��^CzE=���Xs@A}�����@|D�>Z�z��"�}��r��x�:9�:���	��h�D��ُX�Թ*j�Ԛ�#J''�-�&�S���b�޶[ ��&Jx��;�cW�3�zM�H��o���iM����J!�7
�z떠*U?�������I�ԐTt^���$9A��ò*�ژ�Y��Tjc���n�:#��au$£qiH�����2�sfl��I�E/!T��-�fn<�����8ZL�q�]:��N&� b��솞��������6�l3�U��.	����z��@#����Rs�Uӓ����4�K*��u�-���ǎ�5�J$�q�XS/�fwr��5Ӟ�	�
�A�(0��JC]!V)�H#\	#��S�c�7J�3D@x��C?].-H(��bw��d��/9� -��Uӵ��/�n]j�̒�/�:p�ZZ?����R�g���Ƞ-��U�~]=�sk�L/�r�=�3���O�Q��Z�@"qj��i��Nb�rN~7j�$M�~�n�l6��+CҶ�x��Р��.1�Jc�qls�߾,fZ��kq9�j{z�it�wXo���Y��XJ!��e�Պ��Hz��X{��/����+_1���ԓ �d��0���h)_�8hܩ��2��+�����OT��Y��]�����-�D�����;`3���-�L�Lh^�S����0�չe-'������E��PYL檻�(e,op�G��ڮQ#���/�?�Q���Yڈw4�H���z����S�m��[Bf���߱�b�������}1}��7�>�.����4��W>a��Г��0
���R	�t�h:�*Ug���	/Vˉ8�0�HG�f���o�o_�|F��
�Ms�V��n�Q�ھƼ��sc�q��R��6cF�[�&���������6�%"��j�q*�fM�����s��d3G1��W�������nv��E�p��@�p�I�.�˜�O�쯞?��R���������{����|wPJ���L̙�ɾ�^�B��5�l���'��r�;������}JCWC�[��]6��ឈ� >�ͻ;Z��    IEND�B`�