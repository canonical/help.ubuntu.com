<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Mittenklick</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> › <a class="trail" href="mouse.html#tips" title="Tips">Tips</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> › <a class="trail" href="mouse.html#tips" title="Tips">Tips</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="tips.html" title="Tips och tricks">Tips och tricks</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Mittenklick</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Många möss och styrplattor har en musknapp mellan vänster och höger knapp. På en mus med rullningshjul kan du i regel trycka ner själva hjulet för att mittenklicka. Om du inte har en mittenknapp kan du trycka ner vänster och höger musknappar samtidigt för att mittenklicka. Om du ändå inte kan mittenklicka på det här sättet kan du prova att följa <span class="link"><a href="https://wiki.ubuntu.com/X/Quirks#A2-button_Mice" title="https://wiki.ubuntu.com/X/Quirks#A2-button_Mice">dessa instruktioner</a></span>.</p>
<p class="p">På styrplattor som har stöd för flerfingergester kan du peka med tre fingrar samtidigt för att mittenklicka. Du måste <span class="link"><a href="mouse-touchpad-click.html" title="Klicka, dra, eller rulla med styrplattan">aktivera pek-klick</a></span> i styrplatteinställningarna för att det här ska fungera.</p>
<p class="p">Många program använder mittenklick för avancerade klick-kommandon.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list">
<p class="p">Ett vanligt klick-kommando är att klistra in markerad text. (Detta kallas ibland primär markeringsklistring.) Markera texten du vill klistra in, och gå sedan dit du vill klistra in den och mittenklicka. Den markerade texten klistras in vid muspekaren.</p>
<p class="p">Att klistra in text med din mittenknapp sker helt separat från det vanliga klippbordet. Att markera text kopierar den inte till ditt klippbord. Den här snabba metoden för att klistra in fungerar bara med musens mittenknapp.</p>
</li>
<li class="list"><p class="p">I rullningslister och reglage flyttar ett enkelklick i den tomma ytan ett visst avstånd (till exempel en sida) i den riktningen du klickade i. Du kan också mittenklicka i det tomma området för att flytta till just den plats du klickade på.</p></li>
<li class="list"><p class="p">Du kan snabbt öppna ett nytt fönster för ett program med ett mittenklick. Mittenklicka på programmets ikon, antingen i <span class="gui">Startaren</span> till vänster, eller i <span class="gui">Dash</span>.</p></li>
<li class="list"><p class="p">De flesta webbläsare låter dig snabbt öppna länkar i flikar med musens mittenknapp. Klicka på någon länk med din mittenknapp, så öppnas den i en ny flik. Var bara försiktig om du klickar på länken i webbläsaren <span class="app">Firefox</span>. I <span class="app">Firefox</span>, om du mittenklickar någon annanstans än på en länk kommer den försöka läsa den markerade texten som en URL, som om du använda mittenklick för att klistra in den i platsraden och tryckte <span class="key"><kbd>Retur</kbd></span>.</p></li>
<li class="list"><p class="p">I filhanteraren har mittenklick två roller. Om du mittenklickar på en mapp kommer den öppnas i en ny flik. Detta härmar beteendet i vissa populära webbläsare. Om du mittenklickar på en fil kommer den öppnas, precis som om du dubbelklickade.</p></li>
</ul></div></div></div>
<p class="p">Vissa specialiserade program låter dig använda mittenknappen för andra funktioner. Sök i ditt programs hjälpdokument för <span class="em">mittenklick</span> eller <span class="em">musens mittknapp</span>.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="mouse.html#tips" title="Tips">Mustips</a></li>
<li class="links ">
<a href="tips.html" title="Tips och tricks">Tips och tricks</a><span class="desc"> — <span class="link"><a href="tips-specialchars.html" title="Skriv speciella tecken">Speciella tecken</a></span>, <span class="link"><a href="mouse-middleclick.html" title="Mittenklick">mittenklick</a></span>…</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
