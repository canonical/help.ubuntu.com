<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Starta program</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="getting-started.html" title="Komma igång">Börja med GNOME</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks"><a class="nextlinks-next" href="gs-switch-tasks.html" title="Växla uppgifter">Nästa</a></div>
<div class="hgroup"><h1 class="title"><span class="title">Starta program</span></h1></div>
<div class="region">
<div class="contents"><div class="ui-tile ">
<a href="figures/gnome-launching-applications.webm" class="ui-overlay"><span class="ui-tile-img" style="width: 812px; height: 452px;"><img src="gs-thumb-launching-apps.svg" width="812" height="452"></span></a><div class="ui-overlay"><div class="inner">
<a href="#" class="ui-overlay-close" title="Stäng">⨯</a><div class="contents"><div class="media media-video"><div class="inner">
<video src="figures/gnome-launching-applications.webm" preload="auto" controls="controls" class="media media-block" height="394" width="700" data-play-label="Spela upp" data-pause-label="Paus"></video><div class="media-ttml">
<div class="media-ttml-node media-ttml-div" data-ttml-begin="1" data-ttml-end="5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="1" data-ttml-end="5">Starta program</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="5" data-ttml-end="7.5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="5" data-ttml-end="7.5">Flytta din musmarkör till <span class="gui">Aktivitetshörnet</span> längst upp till vänster på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="7.5" data-ttml-end="9.5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="7.5" data-ttml-end="9.5">Klicka på ikonen <span class="gui">Visa program</span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="9.5" data-ttml-end="11"><div class="media-ttml-node media-ttml-p" data-ttml-begin="9.5" data-ttml-end="11">Klicka på programmet som du vill köra, till exempel, Hjälp.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="12" data-ttml-end="21"><div class="media-ttml-node media-ttml-p" data-ttml-begin="12" data-ttml-end="21">Alternativt, använd tangentbordet för att öppna <span class="gui">Aktivitetsöversikt</span> genom att trycka på <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="22" data-ttml-end="29"><div class="media-ttml-node media-ttml-p" data-ttml-begin="22" data-ttml-end="29">Börja skriva namnet på det program du vill starta.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="30" data-ttml-end="33"><div class="media-ttml-node media-ttml-p" data-ttml-begin="30" data-ttml-end="33">Tryck på <span class="key"><kbd>Retur</kbd></span> för att starta programmet.</div></div>
</div>
</div></div></div>
</div></div>
</div></div>
<div id="launch-apps-mouse" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Starta program med musen</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Flytta din musmarkör till <span class="gui">Aktivitetshörnet</span> längst upp till vänster på skärmen för att visa <span class="gui">Aktivitetsöversikt</span>.</p></li>
<li class="steps"><p class="p">Klicka på ikonen <span class="gui">Visa program</span> som visas i botten av panelen i vänstersidan på skärmen.</p></li>
<li class="steps"><p class="p">En lista av program visas. Klicka på programmet som du vill köra, till exempel Hjälp.</p></li>
</ol></div></div></div></div></div>
</div></div>
<div id="launch-app-keyboard" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Starta program med tangentbordet</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna <span class="gui">Aktivitetsöversikt</span> genom att trycka på <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>.</p></li>
<li class="steps"><p class="p">Börja skriv namnet på programmet som du vill starta. Sökningen efter programmet påbörjas omedelbart.</p></li>
<li class="steps"><p class="p">När programmets ikon visas och är markerad, tryck på <span class="key"><kbd>Retur</kbd></span> för att starta programmet.</p></li>
</ol></div></div></div></div></div>
</div></div>
<div class="links nextlinks"><a class="nextlinks-next" href="gs-switch-tasks.html" title="Växla uppgifter">Nästa</a></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="getting-started.html" title="Komma igång">Börja med GNOME</a><span class="desc"> — Är GNOME nytt för dig? Lär dig hur du använder det.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-apps-open.html" title="Starta program">Starta program</a><span class="desc"> — Starta program från översiktsvyn <span class="gui">Aktiviteter</span>.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
