<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Användarkonton</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 23.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Användarkonton</span></h1></div>
<div class="region">
<div class="contents pagewide"><p class="p">Varje person som använder datorn bör ha ett eget användarkonto. Detta låter dem ha sina filer separat från dina och att välja sina egna inställningar. Det är också säkrare. Du kan bara nå ett annat användarkonto om du vet dess lösenord.</p></div>
<section id="manage"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Hantera användarkonton</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="user-add.html.sv" title="Lägg till ett nytt användarkonto"><span class="title">Lägg till ett nytt användarkonto</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till nya användare så att andra personer kan logga in på datorn.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-autologin.html.sv" title="Logga in automatiskt"><span class="title">Logga in automatiskt</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in automatisk inloggning när du startar din dator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="parental-controls.html.sv" title="Lägg till föräldrakontroller"><span class="title">Lägg till föräldrakontroller</span><span class="linkdiv-dash"> — </span><span class="desc">Konfigurera föräldrakontroller för användare på systemet.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="user-delete.html.sv" title="Ta bort ett användarkonto"><span class="title">Ta bort ett användarkonto</span><span class="linkdiv-dash"> — </span><span class="desc">Ta bort användare som inte längre använder din dator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-changepicture.html.sv" title="Ändra ditt foto på inloggningsskärmen"><span class="title">Ändra ditt foto på inloggningsskärmen</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till ditt foto till inloggnings- och användarskärmarna.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="passwords"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Lösenord</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs"><div class="linkdiv "><a class="linkdiv" href="user-changepassword.html.sv" title="Välj ditt lösenord"><span class="title">Välj ditt lösenord</span><span class="linkdiv-dash"> — </span><span class="desc">Håll ditt konto säkert genom att ändra ditt lösenord ofta i dina kontoinställningar.</span></a></div></div>
<div class="links-divs"><div class="linkdiv "><a class="linkdiv" href="user-goodpassword.html.sv" title="Välj ett säkert lösenord"><span class="title">Välj ett säkert lösenord</span><span class="linkdiv-dash"> — </span><span class="desc">Använd längre och mer komplicerade lösenord.</span></a></div></div>
</div></div></div></div></div></div>
</div></section><section id="privileges"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Användarbehörigheter</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="user-admin-explain.html.sv" title="Hur fungerar administratörsbehörighet?"><span class="title">Hur fungerar administratörsbehörighet?</span><span class="linkdiv-dash"> — </span><span class="desc">Du behöver administratörsbehörighet för att ändra viktiga delar i ditt system.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-admin-problems.html.sv" title="Problem som orsakas av administratörsbegränsningar"><span class="title">Problem som orsakas av administratörsbegränsningar</span><span class="linkdiv-dash"> — </span><span class="desc">Vissa saker, som att installera program, kan du endast göra om du har administratörsbehörighet.</span></a></div>
</div>
<div class="links-divs"><div class="linkdiv "><a class="linkdiv" href="user-admin-change.html.sv" title="Ändra vem som har administratörsbehörighet"><span class="title">Ändra vem som har administratörsbehörighet</span><span class="linkdiv-dash"> — </span><span class="desc">Du kan tillåta användare att göra ändringar för systemet genom att ge dem administratörsbehörighet.</span></a></div></div>
</div></div></div></div></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — Få GNOME att arbeta för dig, från hårdvarukontroll till sekretessinställningar.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
