<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="500" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-go-online2.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns1:collect="always" id="linearGradient14901">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop14903"/>
      <ns0:stop style="stop-color:#000000;stop-opacity:0;" offset="1" id="stop14905"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2">
      <ns0:stop id="stop3964-5-0-1-9-6-6" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68893" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:linearGradient id="linearGradient6868-5-7-5-4-3" ns1:collect="always">
      <ns0:stop id="stop6870-84-7-0-1-8" offset="0" style="stop-color: rgb(0, 0, 0); stop-opacity: 1;"/>
      <ns0:stop id="stop6872-0-5-0-7-1" offset="1" style="stop-color: rgb(0, 0, 0); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68891" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68897" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68895" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68901" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68899" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68905" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68903" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68909" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68907" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68913" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68911" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68917" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68915" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68921" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68919" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68925" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3" id="radialGradient68923" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" r="19.18985"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath56767">
      <ns0:path ns2:nodetypes="ccccc" ns1:connector-curvature="0" id="path56769" d="m 228.45991,29.202459 833.57379,0 0,290.286071 c -330.23641,0 -408.68316,175.76954 -833.57379,175.76954 z" style="color:#000000;fill:#babdb6;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath14882">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:8.72566223;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path14884" ns2:cx="2246" ns2:cy="390" ns2:rx="482" ns2:ry="482" d="m 2728,390 a 482,482 0 1 1 -964,0 482,482 0 1 1 964,0 z" transform="matrix(0.35527386,0,0,0.35527386,119.03054,9.4159878)"/>
    </ns0:clipPath>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient14901" id="linearGradient14907" x1="532.43353" y1="187.53497" x2="532.43353" y2="314.62036" gradientUnits="userSpaceOnUse"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-2-7-1">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-4-6-6" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-1-4-3">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-5-5" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-3-9">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-5-4" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25942">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25944" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25946">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25948" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25950">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25952" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-9-6-0">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-1-6-2" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-6-4-2-8">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-19-7-4" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-8-2-8-7-5">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-9-2-7-6-1" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25960">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25962" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25964">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25966" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25968">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25970" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25972">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25974" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25976">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25978" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25980">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25982" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25984">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25986" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25988">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25990" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25992">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25994" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25996">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect25998" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath26000">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect26002" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath26004">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect26006" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath24971-0" clipPathUnits="userSpaceOnUse">
      <ns0:rect y="-354.29291" x="624" height="93" width="276" id="rect24973-5" style="color:#000000;fill:none;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-2-7">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-4-6" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-1-4">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-5" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-3">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-5" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-1-7">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-9-9);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-5-6" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-5-5" id="radialGradient12116-6-2-9-3-0-9-9" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-5-5">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-4-1"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-8-15"/>
    </ns0:linearGradient>
    <ns0:clipPath id="clipPath4201-6-8-5-59">
      <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="path4203-1-2-5-0" ns1:connector-curvature="0" d="m 101,177 0,5 2,0 0,2 1,0 0,-4 7,0 0,4 1,0 0,-2 2,0 0,-5 -13,0 z"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-9-6">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6281-3-1-6" y="220.75" x="26.85" height="6.3750005" width="3.8250003"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-6-4-2">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6267-6-9-19-7" y="221.32954" x="26.96591" height="5.21591" width="2.8977277"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-8-2-8-7">
      <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect6261-4-9-2-7-6" y="221.50153" x="26.998718" height="4.8734746" width="1.8762827"/>
    </ns0:clipPath>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-3-7">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-75-13);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-6-5" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-7-2" id="radialGradient12116-6-2-9-3-0-75-13" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-7-2">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-8-92"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-04-00"/>
    </ns0:linearGradient>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-0-0">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-7-75);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-3-8" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-9-1" id="radialGradient12116-6-2-9-3-0-7-75" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-9-1">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-3-4"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-0-50"/>
    </ns0:linearGradient>
    <ns0:mask maskUnits="userSpaceOnUse" id="mask12112-0-6-5-3-8-4">
      <ns0:rect style="fill:url(#radialGradient12116-6-2-9-3-0-3);fill-opacity:1;stroke:none" id="rect12114-2-9-0-8-2-0" width="221" height="16" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-77" id="radialGradient12116-6-2-9-3-0-3" gradientUnits="userSpaceOnUse" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" cx="128.5" cy="442" fx="128.5" fy="442" r="110.5"/>
    <ns0:linearGradient ns1:collect="always" id="linearGradient12104-5-1-5-6-8-77">
      <ns0:stop style="stop-color:#cccccc;stop-opacity:1;" offset="0" id="stop12106-3-0-0-5-2-87"/>
      <ns0:stop style="stop-color:#cccccc;stop-opacity:0;" offset="1" id="stop12108-4-0-4-9-5-7"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" id="linearGradient14901-1">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop14903-7"/>
      <ns0:stop style="stop-color:#000000;stop-opacity:0;" offset="1" id="stop14905-2"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(0.75098334,0,0,0.75098334,-170.84871,-42.430559)" y2="314.62036" x2="532.43353" y1="187.53497" x1="532.43353" gradientUnits="userSpaceOnUse" id="linearGradient27012" ns4:href="#linearGradient14901-1" ns1:collect="always"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-9">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9-8" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9-6" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6-7" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-6-1">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-3-1" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-33-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-6-5" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-6-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-4-9" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath32041">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect32043" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath32045">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect32047" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-6-8-25-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-4-9-24-2" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-6-1-4-5">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-3-0-3-5" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-33-6-5-1-3">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-6-9-1-4-8" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-6-8-2-1-6-6">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-4-9-2-0-9-0" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:filter color-interpolation-filters="sRGB" ns1:collect="always" x="-0.10291173" width="1.2058235" y="-0.065432459" height="1.1308649" id="filter5601">
      <ns0:feGaussianBlur ns1:collect="always" stdDeviation="0.610872" id="feGaussianBlur5603"/>
    </ns0:filter>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-6" id="linearGradient48287" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient id="linearGradient5716-6">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-7"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-7"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716-6" id="linearGradient48289" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:linearGradient id="linearGradient33938">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop33940"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop33942"/>
    </ns0:linearGradient>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient33948" ns4:href="#linearGradient5716-6" ns1:collect="always"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-7">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9-2" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4-0">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9-2" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2-5">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6-2" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="-204.5363" ns1:cy="342.43398" ns1:document-units="px" ns1:current-layer="g26899" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="5120" ns1:window-height="1376" ns1:window-x="0" ns1:window-y="27" ns1:window-maximized="1" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="656" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-540)">
    <ns0:g id="g27126" transform="translate(9,-167.29113)">
      <ns0:g id="g15031" transform="translate(-51,24.637831)">
        <ns0:path transform="translate(2,453.36217)" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" ns2:ry="17" ns2:rx="17" ns2:cy="278" ns2:cx="120" id="path15033" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
        <ns0:text id="text15035" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan15037" ns2:role="line" style="font-size:14px;line-height:1.25">1</ns0:tspan></ns0:text>
      </ns0:g>
      <ns0:g clip-path="none" transform="matrix(0.7432991,0,0,0.7432991,3.7849383,392.29986)" id="g26899">
        <ns0:path style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2.93785119;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 659.42842,512.06341 c -0.7509,0 -1.48468,0.26524 -2.06007,0.84084 l -23.88003,23.88003 -308.21205,0 c -6.5103,0 -11.77184,5.26154 -11.77184,11.77184 l 0,164.46945 427.444,0 0,-164.46945 c 0,-6.5102 -5.2196,-11.77184 -11.7298,-11.77184 l -43.85012,0 -23.88002,-23.88003 c -0.5755,-0.5754 -1.30917,-0.84084 -2.06007,-0.84084 z m -345.92399,348.95104 0,132.47526 c 0,6.51019 5.26154,11.77189 11.77184,11.77189 l 403.94236,0 c 6.5102,0 11.7298,-5.2617 11.7298,-11.77189 l 0,-132.47526 z" id="rect41123-4" ns1:connector-curvature="0" ns2:nodetypes="sccssccssccscsssscc"/>
        <ns0:g transform="matrix(3.7117385,0,0,3.7117385,441.75165,732.88835)" ns1:label="#g5607" id="default-pointer-c" style="display:inline">
          <ns0:path ns2:nodetypes="cccccccc" id="path5567" d="m 27.135224,2.8483222 0,16.4402338 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 27.135224,2.8483222 z" style="opacity:0.6;color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;filter:url(#filter5601);enable-background:accumulate" ns1:connector-curvature="0"/>
          <ns0:path style="color:#000000;fill:url(#linearGradient48287);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path5565" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
          <ns0:path ns2:nodetypes="cccccccc" id="path6242" d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" style="color:#000000;fill:url(#linearGradient33948);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
        </ns0:g>
        <ns0:g id="g15062" transform="matrix(1.3453534,0,0,1.3453534,332.63788,598.67052)" style="fill:#000000;fill-opacity:1;display:inline">
          <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" id="g15066" transform="translate(-81,-317)" ns1:label="status">
            <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" id="g15068" transform="translate(0,40)">
              <ns0:rect style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="2.9722719" height="2" ry="0.5625" rx="0.5625" id="rect15070" y="284" x="81"/>
              <ns0:rect style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="3.0164659" height="2" ry="0.5625" rx="0.5625" id="rect15072" y="284" x="93.983536"/>
            </ns0:g>
            <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" id="g15074" transform="matrix(0.70710678,-0.70710679,0.70710679,0.70710678,-175.45794,186.40707)">
              <ns0:rect width="2.9722719" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ry="0.5625" height="2" rx="0.5625" id="rect15076" y="284" x="81"/>
              <ns0:rect width="3.0164659" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ry="0.5625" height="2" rx="0.5625" id="rect15078" y="284" x="93.983536"/>
            </ns0:g>
            <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" id="g15080" transform="matrix(0,-1,1,0,-196,414)">
              <ns0:rect style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="2.9722719" height="2" ry="0.5625" rx="0.5625" id="rect15082" y="284" x="81"/>
              <ns0:rect style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="3.0164659" height="2" ry="0.5625" rx="0.5625" id="rect15084" y="284" x="93.983536"/>
            </ns0:g>
            <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" id="g15086" transform="matrix(-0.70710679,-0.70710678,0.70710678,-0.70710679,-49.592928,589.45794)">
              <ns0:rect width="2.9722719" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ry="0.5625" height="2" rx="0.5625" id="rect15088" y="284" x="81"/>
              <ns0:rect width="3.0164659" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ry="0.5625" height="2" rx="0.5625" id="rect15090" y="284" x="93.983536"/>
            </ns0:g>
            <ns0:path style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2.16944861;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans" id="path15092" d="m 89.034905,320.9942 c -2.171787,0 -3.946856,1.77507 -3.946856,3.94686 0,2.17178 1.775069,3.97566 3.946856,3.97566 2.171787,0 3.975664,-1.80388 3.975664,-3.97566 0,-2.17179 -1.803877,-3.94686 -3.975664,-3.94686 z m 0,2.01664 c 1.090904,0 1.959023,0.83931 1.959023,1.93022 0,1.0909 -0.868119,1.95902 -1.959023,1.95902 -1.090904,0 -1.930214,-0.86812 -1.930214,-1.95902 0,-1.09091 0.83931,-1.93022 1.930214,-1.93022 z" ns1:connector-curvature="0"/>
          </ns0:g>
          <ns0:g id="g15094" transform="translate(-81,-317)" ns1:label="devices" style="fill:#ffffff;fill-opacity:1"/>
          <ns0:g id="g15096" transform="translate(-81,-317)" ns1:label="apps" style="fill:#ffffff;fill-opacity:1"/>
          <ns0:g id="g15098" transform="translate(-81,-317)" ns1:label="actions" style="fill:#ffffff;fill-opacity:1"/>
          <ns0:g id="g15100" transform="translate(-81,-317)" ns1:label="places" style="fill:#ffffff;fill-opacity:1"/>
          <ns0:g id="g15102" transform="translate(-81,-317)" ns1:label="mimetypes" style="fill:#ffffff;fill-opacity:1"/>
          <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" id="g15104" transform="translate(-81,-317)" ns1:label="emblems"/>
          <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" id="g15106" transform="translate(-81,-317)" ns1:label="categories"/>
        </ns0:g>
        <ns0:rect ry="1.7873727" rx="1.8594906" y="-720.68964" x="607.55249" height="345.7753" width="3.7617662" id="rect15756" style="color:#000000;fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1.32587242;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(0,1,-1,0,0,0)"/>
        <ns0:path ns2:type="arc" style="fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1;stroke-opacity:1;display:inline" id="path15762" ns2:cx="853.0816" ns2:cy="116.95945" ns2:rx="3.6702957" ns2:ry="3.6702957" d="m 856.7519,116.95945 c 0,2.02705 -1.64325,3.6703 -3.6703,3.6703 -2.02704,0 -3.67029,-1.64325 -3.67029,-3.6703 0,-2.02705 1.64325,-3.6703 3.67029,-3.6703 2.02705,0 3.6703,1.64325 3.6703,3.6703 z" transform="matrix(0,2.6014918,-2.6014918,0,910.14466,-1609.8514)"/>
        <ns0:rect transform="matrix(0,1,-1,0,0,0)" style="color:#000000;fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1.32587242;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect59830" width="3.7617662" height="345.7753" x="569.88251" y="-720.68964" rx="1.8594906" ry="1.7873727"/>
        <ns0:path transform="matrix(0,2.6014918,-2.6014918,0,955.88668,-1647.5213)" d="m 856.7519,116.95945 c 0,2.02705 -1.64325,3.6703 -3.6703,3.6703 -2.02704,0 -3.67029,-1.64325 -3.67029,-3.6703 0,-2.02705 1.64325,-3.6703 3.67029,-3.6703 2.02705,0 3.6703,1.64325 3.6703,3.6703 z" ns2:ry="3.6702957" ns2:rx="3.6702957" ns2:cy="116.95945" ns2:cx="853.0816" id="path59832" style="fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1;stroke-opacity:1;display:inline" ns2:type="arc"/>
        <ns0:g style="fill:#ffffff;fill-opacity:1;display:inline" ns1:label="audio-speakers" transform="matrix(1.3453534,0,0,1.3453534,308.37527,269.05896)" id="g5525-4-0">
          <ns0:path style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" d="m 27.433982,218 -3.84375,4.03125 -3.5625,0 0,6.125 3.5625,0 3.9375,3.84375 0.5,-0.0312 0,-13.9375 z" id="path5533-7" ns1:connector-curvature="0" ns2:nodetypes="ccccccccc"/>
          <ns0:path style="fill:none;stroke:#ffffff;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" d="m 30.939342,221 2,-2" id="path8311" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
          <ns0:path ns1:connector-curvature="0" id="path9081" d="m 30.939342,229 2,2" style="fill:none;stroke:#ffffff;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns2:nodetypes="cc"/>
          <ns0:path style="color:#000000;fill:none;stroke:#ffffff;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="m 31.939342,225.0202 3.03125,0" id="path9083" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
          <ns0:rect style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect9102" width="1.0000017" height="1" x="29.93936" y="221"/>
          <ns0:rect y="228" x="29.93936" height="1" width="1.0000017" id="rect9104" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
        </ns0:g>
        <ns0:rect style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect59873" width="429.16772" height="44.396664" x="312.41132" y="668.62891" rx="0" ry="0"/>
        <ns0:text id="text32132" y="698.00366" x="366.59216" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" xml:space="preserve"><ns0:tspan y="698.00366" x="366.59216" id="tspan32134" ns2:role="line" style="font-size:20.56496048px;line-height:1.25">Trådlöst nätverk</ns0:tspan></ns0:text>
        <ns0:g style="display:inline" transform="matrix(1.3453534,0,0,1.3453534,274.74144,415.70247)" id="g3944" ns1:label="network-wireless-signal-good">
          <ns0:path clip-path="url(#clipPath6279-6-1)" ns2:type="arc" style="fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path3743" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" transform="matrix(0,-0.784314,0.784314,0,-128.137,227.059)" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
          <ns0:path clip-path="url(#clipPath6265-33-4)" transform="matrix(0,-1.72549,1.72549,0,-338.902,250.529)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3745-5" style="fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" ns2:type="arc" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
          <ns0:rect transform="matrix(0,-1,1,0,0,0)" ns1:label="audio-volume-high" y="40" x="-212" height="16" width="16" id="rect3749" style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible"/>
          <ns0:path transform="matrix(1.5,0,0,1.5,5.5,-105)" d="m 29,209 c 0,0.55228 -0.447715,1 -1,1 -0.552285,0 -1,-0.44772 -1,-1 0,-0.55228 0.447715,-1 1,-1 0.552285,0 1,0.44772 1,1 z" ns2:ry="1" ns2:rx="1" ns2:cy="209" ns2:cx="28" id="path3751" style="fill:#000000;fill-opacity:1;stroke:none;display:inline" ns2:type="arc"/>
          <ns0:path ns2:end="7.0685835" ns2:start="5.4977871" ns2:open="true" transform="matrix(0,-2.66667,2.66667,0,-549.666,274)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path2937-7" style="opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" ns2:type="arc" clip-path="url(#clipPath6259-6-8-25-4)"/>
        </ns0:g>
        <ns0:text xml:space="preserve" style="color:#000000;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-indent:0;text-align:end;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:end;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="698.89441" y="698.00366" id="text59875"><ns0:tspan ns2:role="line" id="tspan59877" x="698.89441" y="698.00366" style="font-size:20.56496048px;line-height:1.25">hemmanätverk</ns0:tspan></ns0:text>
        <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="rect12003" d="m 726.44385,688.97738 -5.04507,5.04508 -5.04509,-5.04508 z" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
        <ns0:text xml:space="preserve" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="331.61298" y="753.16315" id="text59897"><ns0:tspan ns2:role="line" id="tspan59899" x="331.61298" y="753.16315" style="font-size:20.56496048px;line-height:1.25">Välj nätverk</ns0:tspan></ns0:text>
        <ns0:text id="text59901" y="796.2146" x="331.61298" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" xml:space="preserve"><ns0:tspan y="796.2146" x="331.61298" id="tspan59903" ns2:role="line" style="font-size:20.56496048px;line-height:1.25">Stäng av</ns0:tspan></ns0:text>
        <ns0:text xml:space="preserve" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="331.61298" y="839.26605" id="text59905"><ns0:tspan ns2:role="line" id="tspan59907" x="331.61298" y="839.26605" style="font-size:20.56496048px;line-height:1.25">Inställningar för trådlösa nätverk</ns0:tspan></ns0:text>
        <ns0:g style="display:inline" ns1:label="audio-volume-medium" transform="matrix(1.3453534,0,0,1.3453534,590.89949,182.95633)" id="g5525">
          <ns0:path ns1:connector-curvature="0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none" d="m 20,222 h 2.484375 L 25.453129,219 26,219.0156 v 11 l -0.475297,8.3e-4 L 22.484375,227 H 20 Z" id="path5533" ns2:nodetypes="ccccccccc"/>
          <ns0:rect ns1:label="audio-volume-high" y="217" x="20" height="16" width="16" id="rect5535" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none"/>
          <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3718-5" style="display:inline;fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:type="arc" clip-path="url(#clipPath6279-7-9-7)"/>
          <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" ns2:type="arc" style="display:inline;fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" id="path3726-1" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" clip-path="url(#clipPath6265-3-4-4-0)"/>
          <ns0:path ns2:end="0.78539819" ns2:start="5.4977871" ns2:open="true" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3728-0" style="display:inline;opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:type="arc" clip-path="url(#clipPath6259-8-81-2-5)"/>
        </ns0:g>
        <ns0:g style="display:inline" id="g4692-3" ns1:label="system-shutdown" transform="matrix(1.3453534,0,0,1.3453534,591.45102,-450.08783)">
          <ns0:rect width="16" height="16" rx="0.14408804" ry="0.15129246" x="40" y="688" id="rect10837-3-0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none;enable-background:new"/>
          <ns0:path ns2:type="arc" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" id="path3869-2" ns2:cx="48" ns2:cy="696" ns2:rx="7" ns2:ry="7" d="m 51.52343,689.95141 a 7,7 0 0 1 3.233191,7.87837 7,7 0 0 1 -6.766907,5.17021 7,7 0 0 1 -6.751683,-5.19008 7,7 0 0 1 3.25633,-7.86883" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" ns2:start="5.239857" ns2:end="4.1878597" ns2:open="true"/>
          <ns0:path ns1:connector-curvature="0" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" d="m 48,689 v 5" id="path4710" ns2:nodetypes="cc"/>
        </ns0:g>
        <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:4.03606033;marker:none;enable-background:accumulate" d="m 685.77004,486.8382 -5.04507,5.04509 -5.04508,-5.04509 z" id="rect12003-0" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
        <ns0:g style="display:inline;enable-background:new" ns1:label="network-wired" id="g8415" transform="matrix(1.3453534,0,0,1.3453534,262.633,236.77047)">
          <ns0:rect y="177" x="241.0002" height="16" width="16" id="rect8417" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none"/>
          <ns0:rect ry="0" y="188" x="241.0002" height="4.9375" width="5.0000014" id="rect8421" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate"/>
          <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate" id="rect8425" width="5.0000014" height="5.0000024" x="251.0002" y="188" ry="0"/>
          <ns0:path style="fill:none;stroke:#1e2224;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" d="M 2.53125,-8.4687501 V -11.5 H 12.5 v 3.0312499" id="path8427" ns1:connector-curvature="0" transform="translate(241.0002,197)" ns2:nodetypes="cccc"/>
          <ns0:path style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" d="M 7.5,-11.5 V -15" id="path9198" ns1:connector-curvature="0" transform="translate(241.0002,197)"/>
          <ns0:rect ry="0" y="178" x="246.0002" height="5.0000024" width="5.0000014" id="rect9200" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate"/>
        </ns0:g>
      </ns0:g>
    </ns0:g>
  </ns0:g>
</ns0:svg>
