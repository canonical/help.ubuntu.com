<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>PHP - Scripting Language</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = "index.html.en";
        } else {
                window.location = href.replace(/\.html.*/, ".html.en");
        }
         return false;
      }
      function browserPreferredLanguage() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = href;
        } else {
                window.location = href.replace(/\.html.*/, ".html");
        }
        return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../18.04" class="trail">Ubuntu 18.04</a> » <a class="trail" href="index.html.sv" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="web-servers.html.sv" title="Webbservrar">Webbservrar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="httpd.html.sv" title="HTTPD - webbservern Apache2">Föregående</a><a class="nextlinks-next" href="squid.html.sv" title="Squid - Proxyserver">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">PHP - Scripting Language</h1></div>
<div class="region">
<div class="contents">
<p class="para">PHP is a general-purpose scripting language suited for Web
      development. PHP scripts can be embedded into HTML. This
      section explains how to install and configure PHP in an Ubuntu
      System with Apache2 and MySQL.</p>
<p class="para"> This section assumes you have installed and configured
      Apache2 Web Server and MySQL Database Server. You can refer to
      the Apache2 and MySQL sections in this document to install and
      configure Apache2 and MySQL respectively.</p>
</div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="php.html.sv#php-installation" title="Installation">Installation</a></li>
<li class="links"><a class="xref" href="php.html.sv#php-configuration" title="Konfiguration">Konfiguration</a></li>
<li class="links"><a class="xref" href="php.html.sv#php-testing" title="Testa">Testa</a></li>
<li class="links"><a class="xref" href="php.html.sv#php-references" title="Referenser">Referenser</a></li>
</ul></div>
<div class="sect2 sect" id="php-installation"><div class="inner">
<div class="hgroup"><h2 class="title">Installation</h2></div>
<div class="region"><div class="contents">
<p class="para">PHP is available in Ubuntu Linux. Unlike python and
      perl, which are installed in the base system, PHP must be added.
      </p>
<div class="steps"><div class="inner"><ul class="steps"><li class="steps">
<p class="para">
      To install PHP and the Apache PHP module you
      can enter the following command at a terminal prompt:

<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install php libapache2-mod-php</span>
</pre></div>
</p>

      <p class="para">You can run PHP scripts at a terminal prompt. To run PHP scripts 
      at a terminal prompt you should install the
      <span class="app application">php-cli</span> package. To install
      <span class="app application">php-cli</span> you can enter the following
      command at a terminal prompt:
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install php-cli</span>
</pre></div>
</p>
      <p class="para">
      You can also execute PHP scripts without installing the Apache PHP
      module. To accomplish this, you should install the
      <span class="app application">php-cgi</span> package. You can run the
      following command at a terminal prompt to install the
      <span class="app application">php-cgi</span> package:
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install php-cgi</span>
</pre></div>
      </p>
      <p class="para">To use <span class="app application">MySQL</span> with PHP you should install
      the <span class="app application">php-mysql</span> package. To install
      <span class="app application">php-mysql</span> you can enter the following
      command at a terminal prompt:
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install php-mysql</span>
</pre></div>
</p>
      <p class="para">Similarly, to use <span class="app application">PostgreSQL</span> with PHP you should install
      the <span class="app application">php-pgsql</span> package. To install
      <span class="app application">php-pgsql</span> you can enter the following
      command at a terminal prompt:
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install php-pgsql</span>
</pre></div>
      </p>
			</li></ul></div></div>
</div></div>
</div></div>
<div class="sect2 sect" id="php-configuration"><div class="inner">
<div class="hgroup"><h2 class="title">Konfiguration</h2></div>
<div class="region"><div class="contents">
<p class="para">
	  If you have installed the
	  <span class="app application">libapache2-mod-php</span> or
	  <span class="app application">php-cgi</span> packages, you can run PHP
	  scripts from your web browser. If you have installed the
	  <span class="app application">php-cli</span> package, you can run PHP
	  scripts at a terminal prompt.
          </p>
<p class="para">
          By default, when <span class="app application">libapache2-mod-php</span>
          is installed, the Apache 2 Web server is configured to run PHP
          scripts. In other words, the PHP module is enabled in the Apache
          Web server when you install the module. Please
          verify if the files
          <span class="file filename">/etc/apache2/mods-enabled/php7.0.conf</span> and
          <span class="file filename">/etc/apache2/mods-enabled/php7.0.load</span>
          exist. If they do not exist, you can enable the module using
          the <span class="cmd command">a2enmod</span> command.
          </p>
<p class="para">Once you have installed the PHP related packages and
	  enabled the Apache PHP module, you should restart the
	  Apache2 Web server to run PHP scripts. You can run the
	  following command at a terminal prompt to restart your web server:
          <div class="screen"><pre class="contents "><span class="cmd command">sudo systemctl restart apache2.service</span> </pre></div>
          </p>
</div></div>
</div></div>
<div class="sect2 sect" id="php-testing"><div class="inner">
<div class="hgroup"><h2 class="title">Testa</h2></div>
<div class="region"><div class="contents">
<p class="para">To verify your installation, you can run the following PHP
          phpinfo script:
          </p>
<div class="code"><pre class="contents ">&lt;?php
  phpinfo();
?&gt;
</pre></div>
<p class="para">
          You can save the content in a file
          <span class="file filename">phpinfo.php</span> and place it
          under the <span class="cmd command">DocumentRoot</span> directory of the
          Apache2 Web server. Pointing your browser to
          <span class="file filename">http://hostname/phpinfo.php</span> will
          display the values of various PHP configuration parameters.
      </p>
</div></div>
</div></div>
<div class="sect2 sect" id="php-references"><div class="inner">
<div class="hgroup"><h2 class="title">Referenser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
            <p class="para">
            For more in depth information see the <a href="http://www.php.net/docs.php" class="ulink" title="http://www.php.net/docs.php">php.net</a> documentation.
            </p> 
          </li>
<li class="list itemizedlist">
            <p class="para">
            There are a plethora of books on PHP.  A good book from O'Reilly is 
            <a href="http://oreilly.com/catalog/0636920043034/" class="ulink" title="http://oreilly.com/catalog/0636920043034/">Learning PHP</a>.
            <a href="http://oreilly.com/catalog/9781565926813/" class="ulink" title="http://oreilly.com/catalog/9781565926813/">PHP Cook Book</a>
            is also good, but has no yet been updated for PHP7.
            </p> 
          </li>
<li class="list itemizedlist">
            <p class="para">
            Also, see the <a href="https://help.ubuntu.com/community/ApacheMySQLPHP" class="ulink" title="https://help.ubuntu.com/community/ApacheMySQLPHP">Apache MySQL PHP Ubuntu Wiki</a> page
            for more information.
            </p> 
          </li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="httpd.html.sv" title="HTTPD - webbservern Apache2">Föregående</a><a class="nextlinks-next" href="squid.html.sv" title="Squid - Proxyserver">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address
          so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>
          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p>
</div>
</div>
</body>
</html>
