<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använd systemsökning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 19.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="getting-started.html.sv" title="Komma igång">Kom igång med GNOME</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<nav class="prevnext pagewide"><div class="inner">
<a href="gs-use-windows-workspaces.html.sv" title="Använda fönster och arbetsytor">Föregående</a><a href="gs-get-online.html.sv" title="Ansluta till nätet">Nästa</a>
</div></nav><div class="hgroup pagewide"><h1 class="title"><span class="title">Använd systemsökning</span></h1></div>
<div class="region">
<div class="contents pagewide">
<div class="media media-image"><div class="inner"><img src="gs-search1.svg" width="100%" class="media media-block" alt=""></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps"><li class="steps">
<p class="p">Öppna översiktsvyn <span class="gui">Aktiviteter</span> genom att klicka på <span class="gui">Aktiviteter</span> högst upp till vänster på skärmen, eller genom att trycka ned knappen <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>. Börja skriva för att söka.</p>
<p class="p">Resultat som matchar det du har skrivit kommer att visas medan du skriver. Det första resultatet är alltid markerat och visas i längst upp.</p>
<p class="p">Tryck på <span class="key"><kbd>Retur</kbd></span> för att växla till det första, markerade resultatet.</p>
</li></ol></div></div></div>
<div class="media media-image"><div class="inner"><img src="gs-search2.svg" width="100%" class="media media-block" alt=""></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps" start="2">
<li class="steps">
<p class="p">Alternativ som kan komma att visas bland sökresultaten inkluderar:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">program som matchar, visas överst bland sökresultaten,</p></li>
<li class="list"><p class="p">matchande inställningar,</p></li>
<li class="list"><p class="p">matchande kontakter,</p></li>
<li class="list"><p class="p">matchande dokument,</p></li>
<li class="list"><p class="p">matchande kalender,</p></li>
<li class="list"><p class="p">matchande kalkylator,</p></li>
<li class="list"><p class="p">matchande programvara,</p></li>
<li class="list"><p class="p">matchande filer,</p></li>
<li class="list"><p class="p">matchande terminal,</p></li>
<li class="list"><p class="p">matchande lösenord och nycklar.</p></li>
</ul></div></div></div>
</li>
<li class="steps">
<p class="p">Bland sökresultaten, klicka på alternativet för att växla till det.</p>
<p class="p">Alternativt, markera ett alternativ genom att använda piltangenterna och tryck på <span class="key"><kbd>Retur</kbd></span>.</p>
</li>
</ol></div></div></div>
</div>
<section id="use-search-inside-applications"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Sök inifrån program</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">Systemsökningen samlar ihop resultat från olika program. Till vänster om sökresultaten kan du se ikoner för de program som tillhandahållit sökresultaten. Klicka på en av ikonerna för att starta om sökningen inifrån programmet som associerats med den ikonen. Eftersom endast de bästa matchningarna visas i <span class="gui">Aktivitetsöversikt</span>, så kan sökning inifrån programmet komma att ge dig bättre sökresultat.</p></div></div>
</div></section><section id="use-search-customize"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Anpassa sökresultat</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="media media-image"><div class="inner"><img src="gs-search-settings.svg" width="100%" class="media media-block" alt=""></div></div>
<div class="note note-important" title="Viktigt">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m12.5 2a9.5 9.5 0 0 0-9.5 9.5 9.5 9.5 0 0 0 9.5 9.5 9.5 9.5 0 0 0 9.5-9.5 9.5 9.5 0 0 0-9.5-9.5zm0 3a1.5 1.5 0 0 1 1.5 1.5v6a1.5 1.5 0 0 1-1.5 1.5 1.5 1.5 0 0 1-1.5-1.5v-6a1.5 1.5 0 0 1 1.5-1.5zm0 10.5a1.5 1.5 0 0 1 1.5 1.5 1.5 1.5 0 0 1-1.5 1.5 1.5 1.5 0 0 1-1.5-1.5 1.5 1.5 0 0 1 1.5-1.5z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Din dator låter dig anpassa vad du vill ska visas bland sökresultaten i <span class="gui">Aktivitetsöversikt</span>. Till exempel så kan du välja om du vill visa resultat för webbplatser, foto eller musik.</p></div></div></div>
</div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">För att anpassa vad som ska visas bland sökresultaten:</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="gui"><a href="shell-introduction.html.sv#yourname" title="shell-introduction#yourname">systemmenyn</a></span> på höger sida av systemraden.</p></li>
<li class="steps"><p class="p">Tryck på inställningsknappen längst ner till vänster i menyn.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Sök</span> i den vänstra panelen.</p></li>
<li class="steps"><p class="p">I listan över sökplatser, klicka på brytaren intill sökplatsen som du vill aktivera eller inaktivera.</p></li>
</ol></div>
</div></div>
</div></div>
</div></section><nav class="prevnext pagewide"><div class="inner">
<a href="gs-use-windows-workspaces.html.sv" title="Använda fönster och arbetsytor">Föregående</a><a href="gs-get-online.html.sv" title="Ansluta till nätet">Nästa</a>
</div></nav><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="getting-started.html.sv" title="Komma igång">Kom igång med GNOME</a><span class="desc"> — Är GNOME nytt för dig? Lär dig hur du använder det.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-apps-open.html.sv" title="Starta program">Starta program</a><span class="desc"> — Starta program från översiktsvyn <span class="gui">Aktiviteter</span>.</span>
</li></ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
