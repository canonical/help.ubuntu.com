<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Redigera en trådlös anslutning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Redigera en trådlös anslutning</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Det här avsnittet beskriver alla alternativ som finns när du redigerar en trådlös nätverksanslutning. För att redigera en anslutning, klicka på <span class="gui">nätverksmenyn</span> i menylisten och välj <span class="gui">Redigera anslutningar</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">De flesta nätverk kommer fungera utmärkt om du lämnar inställningarna orörda, så du behöver antagligen inte ändra något. Många av alternativen här finns till för att ge dig bättre kontroll över mer avancerade nätverk.</p></div></div></div></div>
</div>
<div id="available" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Tillgänglig för alla användare / Anslut automatiskt</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Anslut automatiskt</span></dt>
<dd class="terms">
<p class="p">Kryssa för det här alternativet om du vill att datorn ska försöka ansluta till det här trådlösa nätverket när det finns inom räckhåll.</p>
<p class="p">Om flera nätverk som är inställda för automatisk anslutning finns inom räckhåll kommer datorn ansluta till det som visas överst i fliken <span class="gui">Trådlöst</span> i fönstret <span class="gui">Nätverksanslutningar</span>. Det kommer inte koppla ned från ett tillgängligt nätverk för att ansluta till ett annat som just kom inom räckhåll.</p>
</dd>
<dt class="terms"><span class="gui">Tillgängligt för alla användare</span></dt>
<dd class="terms">
<p class="p">Kryssa för det här om du vill att alla användare på datorn ska kunna komma åt det här trådlösa nätverket. Om nätverket har ett <span class="link"><a href="net-wireless-wepwpa.html" title="Vad betyder WEP och WPA?">WEP-/WPA-lösenord</a></span> och du har kryssat för det här alternativet kommer du bara behöva skriva in lösenordet en gång. Alla andra användare på din dator kommer kunna ansluta till nätverket utan att själva behöva känna till lösenordet.</p>
<p class="p">Om det här är förkryssat behöver du vara en <span class="link"><a href="user-admin-explain.html" title="Hur fungerar administratörsbehörighet?">administratör</a></span> för att ändra inställningar för det här nätverket. Du kan bli ombedd att skriva in ditt administratörslösenord.</p>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div id="wireless" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Trådlöst</span></h2></div>
<div class="region">
<div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">SSID</span></dt>
<dd class="terms"><p class="p">Det här är namnet på det trådlösa nätverk du ansluter till, även kallat <span class="em">Service Set Identifier (SSID)</span>. Ändra inte det här om du inte har ändrat namn på det trådlösa nätverket (genom att till exempel ändra inställningar i din trådlösa router eller basstation).</p></dd>
<dt class="terms"><span class="gui">Läge</span></dt>
<dd class="terms">
<p class="p">Använd det här för att ange om du ansluter till ett <span class="gui">Infrastruktur</span>nätverk (där datorer ansluter trådlöst till en central basstation eller router) eller ett <span class="gui">Ad-hoc</span>-nätverk (där det inte finns någon basstation, och datorerna i nätverket ansluter till varandra). De flesta nätverk är av typen Infrastruktur; du kan dock vilja <span class="link"><a href="net-wireless-adhoc.html" title="Skapa en trådlös surfzon">ställa in ditt eget ad-hoc-nätverk</a></span>.</p>
<p class="p">Om du väljer <span class="gui">Ad-hoc</span> kommer du se två andra alternativ, <span class="gui">Band</span> och <span class="gui">Kanal</span>. Dessa bestämmer vilket trådlöst frekvensband det trådlösa ad-hoc-nätverket ska använda. Vissa datorer kan bara arbeta på vissa band (exempelvis bara <span class="gui">A</span> eller bara <span class="gui">B/G</span>), så du bör välja ett band som alla datorer i ad-hoc-nätverket kan använda. På högtrafikerade platser kan det finnas flera trådlösa nätverk som delar på samma kanal; detta kan sakta ner din anslutning, så du kan också ändra vilken kanal du själv använder.</p>
</dd>
<dt class="terms"><span class="gui">BSSID</span></dt>
<dd class="terms"><p class="p">Det här är <span class="em">Basic Service Set Identifier</span>. SSID:n (se ovan) är namnet på nätverket som det är tänkt att människor ska se; BSSID:n är ett namn som datorn förstår (det är en serie bokstäver och siffror som ska vara unika för det trådlösa nätverket). Om ett <span class="link"><a href="net-wireless-hidden.html" title="Anslut till ett dolt, trådlöst nätverk">nätverl är dolt</a></span> kommer det inte ha en SSID, men det kommer ha en BSSID.</p></dd>
<dt class="terms"><span class="gui">Enhetens MAC-adress</span></dt>
<dd class="terms">
<p class="p">En <span class="link"><a href="net-macaddress.html" title="Vad är en MAC-adress?">MAC-adress</a></span> är en kod som identifierar en nätverkskomponent (till exempel ett trådlöst nätverkskort, ett trådbundet nätverkskort, eller en router). Varje enhet som du kan ansluta till ett nätverk har en unik MAC-adress som tilldelades den vid tillverkning.</p>
<p class="p">Det här alternativet kan användas för att ändra ditt nätverkskorts MAC-adress.</p>
</dd>
<dt class="terms"><span class="gui">Klonad MAC-adress</span></dt>
<dd class="terms"><p class="p">Din nätverkshårdvara (trådlöst kort) kan låtsas ha en annan MAC-adress. Detta kan vara användabart om du har en enhet eller tjänst som bara kommunicerar med en viss MAC-adress (exempelvis ett trådbundet bredbandsmodem). Om du skriver in den MAC-adressen i rutan <span class="gui">klonad MAC-adress</span> kommer enheten/tjänsten tro att din dator har den klonade MAC-adressen istället för den verkliga adressen.</p></dd>
<dt class="terms"><span class="gui">MTU</span></dt>
<dd class="terms"><p class="p">Den här inställningen ändrar <span class="em">maximal överföringsenhet (eng. MTU)</span>, vilket är den största storleken på ett datapaket som kan skickas genom nätverket. När filer skickas genom ett nätverk delas data upp i små paket. Den optimala MTU:n för ditt nätverk kommer bero på hur stor sannolikheten är att paket förloras (på grund av en brusig anslutning) och hur snabb anslutningen är. I allmänhet bör du inte behöva ändra den här inställningen.</p></dd>
</dl></div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless-hidden.html" title="Anslut till ett dolt, trådlöst nätverk">Anslut till ett dolt, trådlöst nätverk</a><span class="desc"> — Klicka på <span class="gui">nätverksmenyn</span> på menylisten och välj <span class="gui">Anslut till dolt trådlöst nätverk</span>.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="security" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Trådlös säkerhet</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Säkerhet</span></dt>
<dd class="terms">
<p class="p">Detta definierar vilken sorts <span class="em">kryptering</span> som ditt trådlösa nätverk använder. Krypterade anslutningar hjälper dig skydda din trådlösa anslutning från avlyssning, så att andra inte kan övervaka dig eller se vilka webbsidor du besöker, osv.</p>
<p class="p">Vissa typer av kryptering är starkare än andra, men kanske inte har lika utbrett stöd av äldre utrustning för trådlösa nätverk. Du kommer i regel behöva skriva in ett lösenord för anslutningen; mer sofistikerade säkerhetstyper kan också kräva ett användarnamn och ett digitalt "certifikat". Se <span class="link"><a href="net-wireless-wepwpa.html" title="Vad betyder WEP och WPA?">Vad betyder WEP och WPA?</a></span> för vidare information om populära typer av trådlös kryptering.</p>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div id="ipv4" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">IPv4-inställningar</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Använd den här fliken för att definiera information som din dators IP-adress och vilka DNS-servrar den bör använda. Ändra <span class="gui">Metod</span> för att se olika sätt att läsa/ändra den informationen.</p>
<p class="p">Följande metoder finns tillgängliga:</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Automatiskt (DHCP)</span></dt>
<dd class="terms"><p class="p">Läs information, som vilken IP-adress och DNS-server som ska användas, från en <span class="em">DHCP-server</span>. En DHCP-server är en dator (eller en annan enhet, som en router) som är ansluten till nätverket som bestämmer vilka nätverksinställningar din dator bör ha - när du först ansluter till nätverket kommer du automatiskt tilldelas lämpliga inställningar. De flesta nätverk använder DHCP.</p></dd>
<dt class="terms"><span class="gui">Endast automatiska (DHCP)-adresser</span></dt>
<dd class="terms"><p class="p">Om du väljer den här inställningen kommer din dator hämta sin IP-adress från en DHCP-server, men du kommer behöva justera övriga detaljer manuellt (som vilken DNS-server du vill använda).</p></dd>
<dt class="terms"><span class="gui">Manuell</span></dt>
<dd class="terms"><p class="p">Välj det här alternativet om du vill definiera alla nätverksinställningar själv, inklusive vilken IP-adress datorn ska använda.</p></dd>
<dt class="terms"><span class="gui">Endast lokal länk</span></dt>
<dd class="terms"><p class="p"><span class="em">Link-Local</span> är ett sätt att ansluta datorer i ett nätverk utan att behöva en DHCP-server eller manuellt definierad IP-adress och annan information. Om du ansluter till ett Link-Local-nätverk kommer datorerna i nätverket själva bestämma vilka IP-adresser som ska användas, och så vidare. Detta är bra om du vill ansluta ett fåtal datorer tillfälligt så att de kan kommunicera med varandra.</p></dd>
<dt class="terms"><span class="gui">Inaktiverad</span></dt>
<dd class="terms"><p class="p">Det här alternativet kommer avaktivera nätverksanslutningen och hindrar dig från att använda den. Observera att <span class="gui">IPv4</span> och <span class="gui">IPv6</span> behandlas som separata anslutningar även om de används av samma nätverkskort. Om en av dem är aktiverad kan du vilja avaktivera den andra.</p></dd>
</dl></div></div></div>
</div></div>
</div></div>
<div id="ipv6" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">IPv6-inställningar</span></h2></div>
<div class="region"><div class="contents"><p class="p">Detta liknar fliken <span class="gui">IPv4</span> förutom att den berör den nyare IPv6-standarden. Moderna nätverk använder IPv6, men IPv4 är i skrivande stund mer populärt.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a><span class="desc"> — <span class="link"><a href="net-wireless-connect.html" title="Anslut till ett trådlöst nätverk">Anslut till trådlöst nätverk</a></span>, <span class="link"><a href="net-wireless-hidden.html" title="Anslut till ett dolt, trådlöst nätverk">Dolda nätverk</a></span>, <span class="link"><a href="net-wireless-edit-connection.html" title="Redigera en trådlös anslutning">Redigera anslutningsinställningar</a></span>, <span class="link"><a href="net-wireless-disconnecting.html" title="Varför kopplar mitt trådlösa nätverk ner hela tiden?">Nedkoppling</a></span>...</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
