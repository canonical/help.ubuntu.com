<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Klicka och flytta muspekaren med det numeriska tangentbordet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="a11y.html" title="Hjälpmedel">Hjälpmedel</a> › <a class="trail" href="a11y.html#mobility" title="Rörelsehinder">Rörelsehinder</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Klicka och flytta muspekaren med det numeriska tangentbordet</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du har svårt att använda en mus eller andra pekdon kan du styra musmarkören via det numeriska tangentbordet på ditt tangentbord. Denna funktion kallas <span class="em">mustangenter</span>.</p>
<p class="p">För att aktivera funktionen mustangenter med hjälp av tangentbordet:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Tryck på <span class="key"><kbd><span class="link"><a href="windows-key.html" title='Vad är "Superknappen"?'>Super</a></span></kbd></span>tangenten för att öppna <span class="gui">Dash</span>.</p></li>
<li class="steps"><p class="p">Skriv <span class="input">Hjälpmedel</span> och tryck <span class="key"><kbd>Retur</kbd></span> för att öppna inställningarna för Hjälpmedel.</p></li>
<li class="steps"><p class="p">Tryck <span class="key"><kbd>Tab</kbd></span> en gång för att välja fliken <span class="gui">Seende</span>.</p></li>
<li class="steps"><p class="p">Tryck <span class="key"><kbd>←</kbd></span> två gånger för att byta till fliken <span class="gui">Peka och klicka</span>.</p></li>
<li class="steps"><p class="p">Tryck <span class="key"><kbd>↓</kbd></span> en gång för att välja växlaren för <span class="gui">Mustangenter</span> och tryck sedan <span class="key"><kbd>Retur</kbd></span> för att slå på dem.</p></li>
<li class="steps"><p class="p">Se till att <span class="key"><kbd>Num Lock</kbd></span> är av. Du kommer nu kunna flytta muspekaren med det numeriska tangentbordet.</p></li>
</ol></div></div></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Ovanstående instruktioner visar det enklaste sättet att aktivera mustangenter genom att bara använda tangentbordet. Välj inställningar för <span class="gui">Hjälpmedel</span> för att se fler åtkomstalternativ.</p></div></div></div></div>
<p class="p"></p>
<p class="p">Det numeriska tangentbordet är en uppsättning sifferknappar på ditt tangentbord, vanligen grupperade i en rektangel. Funktionen mustangenter utgår från tre knappar: den primära, den alternativa och modifiereingsknappen. Nedan följer några exempel på användning av mustangenter:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">Varje siffra på det numeriska tangentbordet (utom 0 och 5) motsvarar en riktning. Till exempel om du trycker på <span class="key"><kbd>8</kbd></span> flyttas markören uppåt och om du trycker på <span class="key"><kbd>2</kbd></span> flyttas den neråt.</p></li>
<li class="list"><p class="p">För att klicka på vald knapp, tryck på <span class="key"><kbd>5</kbd></span>.</p></li>
<li class="list"><p class="p">För att dubbelklicka på vald knapp, tryck på <span class="key"><kbd>5</kbd></span> två gånger eller tryck på <span class="key"><kbd>+</kbd></span> en gång.</p></li>
<li class="list"><p class="p">För att högerklicka, tryck på <span class="key"><kbd>-</kbd></span> för att välja alternativknappen (om den inte redan är vald) och tryck på <span class="key"><kbd>5</kbd></span>.</p></li>
<li class="list"><p class="p">För att mittenklicka, tryck på <span class="key"><kbd>*</kbd></span> för att välja modifieringsknappen (om den inte redan är vald) och tryck på <span class="key"><kbd>5</kbd></span>.</p></li>
<li class="list"><p class="p">För att dra och släppa med hjälp av den primära knappen, tryck på <span class="key"><kbd>/</kbd></span> för att välja den primära knappen (om den inte redan är vald), tryck på <span class="key"><kbd>0</kbd></span> för att trycka ned knappen, dra pekaren dit du önskar, och tryck på <span class="key"><kbd>.</kbd></span> för att släppa knappen.</p></li>
</ul></div></div></div>
<p class="p">
 </p>
<p class="p">Här är en tabell med mustangenter och motsvarande händelser:</p>
<div class="table"><div class="inner"><div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="em">Tangent</span></p></td>
<td><p class="p"><span class="em">Händelse</span></p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>8</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren uppåt</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>2</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren neråt</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>6</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren åt höger</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>4</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren åt vänster</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>7</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren uppåt och åt vänster</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>9</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren uppåt och åt höger</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>3</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren neråt och åt höger</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>1</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Pekaren neråt och åt vänster</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>/</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Välj den primära knappen. På en mus är den primära knappen normalt den vänstra knappen</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>*</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Välj modifieringsknappen. På en mus är modifieringsknappen normalt (om den finns) mellanknappen</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>-</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Välj alternativknappen. På en mus är alternativknappen normalt den högra knappen</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>5</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Klicka på vald knapp</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>+</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Dubbelklicka på vald knapp</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>0</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Tryck på vald knapp</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>,</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Släpp vald knapp</p></td>
</tr>
</table></div></div></div>
<p class="p">
</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om ditt tangentbord saknar ett numeriskt tangentbord (som på en del bärbara datorer), kan du behöva hålla ned funktionstangenten (<span class="key"><kbd class="key-Fn">Fn</kbd></span>) och använda vissa andra tangenter som ett numeriskt tangentbord. Om du använder den här funktionen ofta, kanske du vill köpa ett externt USB-anslutet numeriskt tangentbord.</p></div></div></div></div>
<p class="p">
</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du vill använda det numeriska tangentbordet för att skriva siffror medan mustangenter är aktiverade, slå på <span class="key"><kbd>Num Lock</kbd></span>. Musen kan dock inte styras med det numeriska tangentbordet medan <span class="key"><kbd>Num Lock</kbd></span> är på.</p></div></div></div></div>
<p class="p">
</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">De normala siffertangenterna, i en rad i tangentbordets överkant, kommer inte styra muspekaren. Bara det numeriska tangentbordet kan användas till det här.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="mouse.html" title="Mus">Mus</a><span class="desc"> — <span class="link"><a href="mouse-lefthanded.html" title="Använd din mus med vänster hand">Vänsterhänt</a></span>, <span class="link"><a href="mouse-sensitivity.html" title="Justera hastigheten för musen och styrplattan">hastighet och känslighet</a></span>, <span class="link"><a href="mouse-touchpad-click.html" title="Klicka, dra eller rulla med styrplattan">styrplatteklick och rullning</a></span>…</span>
</li>
<li class="links "><a href="a11y.html#mobility" title="Rörelsehinder">Rörelsehinder</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
