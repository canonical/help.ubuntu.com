<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Tangentbordsnavigation</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="keyboard.html" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="keyboard.html" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="a11y.html" title="Hjälpmedel">Hjälpmedel</a> › <a class="trail" href="a11y.html#mobility" title="Rörelsehinder">Rörelsehinder</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Tangentbordsnavigation</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Denna sida beskriver tangentbordsnavigering för personer som inte kan använda en mus eller annat pekdon eller som vill använda tangentbordet så mycket som möjligt. För snabbtangenter som är användbara för alla användare, se <span class="link"><a href="shell-keyboard-shortcuts.html" title="Användbara tangentbordsgenvägar">Användbara tangentbordsgenvägar</a></span> istället.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du inte kan använda ett pekdon som exempelvis en mus kan du kontrollera musmarkören med hjälp av den numeriska delen på ditt tangentbord. Se <span class="link"><a href="mouse-mousekeys.html" title="Klicka och flytta muspekaren med det numeriska tangentbordet">Klicka och flytta muspekaren med det numeriska tangentbordet</a></span> för detaljer.</p></div></div></div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h2><span class="title">Navigera i användargränssnitt</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="key"><kbd>Tabb</kbd></span> och <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p></td>
<td>
<p class="p">Flytta tangentbordsfokus mellan olika kontroller. <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span> flyttar mellan grupper av kontroller, som exempelvis från en sidopanel till huvudinnehållet. <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span> kan också bryta loss från en kontroll som själv använder <span class="key"><kbd>Tabb</kbd></span>, till exempel ett textområde.</p>
<p class="p">Håll ner <span class="key"><kbd>Skift</kbd></span> för att flytta fokus i omvänd ordning.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Piltangenter</p></td>
<td style="border-top-style: solid;">
<p class="p">Flytta markering mellan objekt i samma kontroll, eller genom en uppsättning relaterade kontroller. Använd piltangenterna för att fokusera på knappar i ett verktygsfält, välj objekt i en list- eller ikonvy, eller välj en radioknapp från en grupp.</p>
<p class="p">I en trädvy, använd vänster och höger piltangent för att fälla ut och ihop objekt med underordnade objekt.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+Piltangenter</span></p></td>
<td style="border-top-style: solid;"><p class="p">I en list- eller ikonvy, flytta tangentbordsfokus till ett annat objekt utan att ändra vilket objekt som är markerat.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Shift</kbd></span>+Piltangenter</span></p></td>
<td style="border-top-style: solid;"><p class="p">I en list- eller ikon-vy, markera alla objekt från och med den för närvarande valda objektet till och med det nyligen fokuserade objektet.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Blanksteg</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Aktivera ett fokuserat objekt som exempelvis en knapp, kryssruta eller listobjekt.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">I en list- eller ikonvy, markera eller avmarkera det fokuserade objektet utan att avmarkera andra objekt.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Alt</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Håll ner <span class="key"><kbd>Alt</kbd></span>-tangenten för att visa <span class="em">snabbtangenter</span>: understrukna bokstäver i menyobjekt, knappar och andra kontroller. Tryck på <span class="key"><kbd>Alt</kbd></span> samt den understrukna bokstaven för att aktivera en kontroll, precis som om du hade klickat på den.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Esc</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Stäng en meny, snabbvalsmeny, växlare eller dialogruta.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>F10</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Öppna den första menyn på menyraden i ett fönster. Använd piltangenterna för att navigera i menyerna.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Shift</kbd></span>+<span class="key"><kbd>F10</kbd></span></span>, eller menytangenten</p></td>
<td style="border-top-style: solid;"><p class="p">Poppa upp snabbvalsmenyn för den aktuella markeringen som om du hade högerklickat.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>F10</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">I filhanteraren, öppna snabbvalsmenyn för den aktuella mappen som om du hade högerklicka på bakgrunden och inte på något objekt.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>PageUp</kbd></span></span> och <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>PageDown</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">I ett gränssnitt med flikar, växla till fliken till vänster eller höger.</p></td>
</tr>
</table></div>
</div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h2><span class="title">Navigera på skrivbordet</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span></p></td>
<td><p class="p"><span class="link"><a href="shell-windows-switching.html" title="Växla mellan fönster">Snabb växling mellan fönster.</a></span> Håll nere <span class="key"><kbd>Shift</kbd></span> för omvänd ordning.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>`</kbd></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p">Växla mellan fönster från samma program, eller från markerat program efter <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span>.</p>
<p class="p">Det här snabbkommandot använder <span class="key"><kbd>`</kbd></span> på amerikanska tangentbord, där tangenten <span class="key"><kbd>`</kbd></span> sitter ovanför <span class="key"><kbd>Tab</kbd></span>. På alla andra tangentbord är kommandot <span class="key"><kbd>Alt</kbd></span> plus vilken tangent som än råkar sitta ovanför <span class="key"><kbd>Tab</kbd></span>.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>piltangenter</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-workspaces-switch.html" title="Växla mellan arbetsytor">Växla mellan arbetsytor.</a></span></p></td>
</tr>
</table></div>
</div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h2><span class="title">Navigera mellan fönster</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F4</kbd></span></span></p></td>
<td><p class="p">Stäng det aktuella fönstret.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><a href="windows-key.html" title='Vad är "Superknappen"?'><kbd>Super</kbd></a></span>+<span class="key"><kbd>↓</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Återställ ett maximerat fönster till dess urspsrungliga storlek.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F7</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Flytta det aktuella fönstret. Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F7</kbd></span></span>, och använd sedan piltangenterna för att flytta fönstret. Tryck <span class="key"><kbd>Retur</kbd></span> för att avsluta flytten, eller <span class="key"><kbd>Esc</kbd></span> för att återgå till den ursprungliga placeringen.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F8</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Ändra storlek på det aktuella fönstret. Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F8</kbd></span></span>, och använd sedan piltangenterna för att ändra fönstrets storlek. Tryck <span class="key"><kbd>Retur</kbd></span> när du är nöjd, eller <span class="key"><kbd>Esc</kbd></span> för att återgå till den ursprungliga storleken.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Shift</kbd></span>+<span class="key"><kbd>piltangenter</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-workspaces-movewindow.html" title="Flytta ett fönster till en annan arbetsyta">Flytta det aktuella fönstret till en annan arbetsyta</a></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><a href="windows-key.html" title='Vad är "Superknappen"?'><kbd>Super</kbd></a></span>+<span class="key"><kbd>↑</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-windows-maximize.html" title="Maximera och avmaximera ett fönster">Maximera</a></span> ett fönster.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><a href="windows-key.html" title='Vad är "Superknappen"?'><kbd>Super</kbd></a></span>+<span class="key"><kbd>←</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Maximera ett fönster vertikalt till vänster på skärmen.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><a href="windows-key.html" title='Vad är "Superknappen"?'><kbd>Super</kbd></a></span>+<span class="key"><kbd>→</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Maximera ett fönster vertikalt till höger på skärmen.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Öppna fönstermenyn, som om du hade högerklickat på namnlisten.</p></td>
</tr>
</table></div>
</div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="a11y.html#mobility" title="Rörelsehinder">Rörelsehinder</a></li>
<li class="links ">
<a href="keyboard.html" title="Tangentbord">Tangentbord</a><span class="desc"> — <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">Indatakällor</a></span>, <span class="link"><a href="keyboard-cursor-blink.html" title="Gör att tangentbordsmarkören blinkar">blinkande markör</a></span>, <span class="link"><a href="windows-key.html" title='Vad är "Superknappen"?'>supertangent</a></span>, <span class="link"><a href="a11y.html#mobility" title="Rörelsehinder">tangentbordsåtkomst</a></span>...</span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-keyboard-shortcuts.html" title="Användbara tangentbordsgenvägar">Användbara tangentbordsgenvägar</a><span class="desc"> — Ta sig runt på skrivbordet med hjälp av tangentbordet.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
