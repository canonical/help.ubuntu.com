<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Visningsinställningar i Filer</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » <a class="trail" href="nautilus-prefs.html" title="Inställningar för filhanterare">Inställningar för filhanterare</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Visningsinställningar i <span class="app">Filer</span></span></h1></div>
<div class="region">
<div class="contents"><p class="p">Du kan ändra standardvyn för nya mappar, hur filer och mappar sorteras, zoomnivån för ikon- och kompaktvyerna, och om filer ska visas i trädvyn bredvid. Välj <span class="guiseq"><span class="gui">Filer</span> ▸ <span class="gui">Inställningar</span></span> i den övre raden medan <span class="app">Filer</span> är öppen och välj fliken <span class="gui">Vyer</span>.</p></div>
<div id="default-view" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Standardvy</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Visa nya mappar med</span></dt>
<dd class="terms"><p class="p">Som standard visas nya mappar i läget ikonvy. Om du föredrar listvyn kan du ställa in det som standard här. Annars kan du välja olika vyer för varje mapp allt eftersom genom att klicka på knappen <span class="gui">Visa objekt som en lista</span> eller <span class="gui">Visa objekt som ikoner</span> i verktygsfältet.</p></dd>
<dt class="terms"><span class="gui">Ordna objekt</span></dt>
<dd class="terms">
<p class="p">Du kan ändra den förvalda sorteringsordningen som används i mappar med den utfällbara listan <span class="gui">Sortera objekt</span> i inställningarna för att sortera efter namn, filstorlek, filtyp, när de senast ändrades, när de senast användas, eller när de togs bort.</p>
<p class="p">Du kan ändra hur <span class="link"><a href="files-sort.html" title="Sortera filer och mappar">filer sorteras</a></span> i en individuell mapp genom att klicka på knappen <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="Visningsalternativ"></span></span> i verktygsfältet och välja <span class="gui">Efter namn</span>, <span class="gui">Efter storlek</span>, <span class="gui">Efter typ</span> eller <span class="gui">Efter ändringsdatum</span>, eller genom att klicka på listkolumnernas rubriker i listvyn. Den här menyn påverkar bara den aktuella mappen.</p>
</dd>
<dt class="terms"><span class="gui">Sortera mappar före filer</span></dt>
<dd class="terms"><p class="p">Som standard visar filhanteraren inte längra alla mappar före filerna. För att se alla mappar ovanför filerna, aktivera det här alternativet.</p></dd>
<dt class="terms"><span class="gui">Visa dolda filer och säkerhetskopior</span></dt>
<dd class="terms">
<p class="p">Filhanteraren visar inte <span class="link"><a href="files-hidden.html" title="Dölj en fil">dolda filer</a></span> och mappar som standard. Du kan alltid visa dolda filer genom att kryssa för det här alternativet.</p>
<p class="p">Du kan också visa dolda filer i ett individuellt fönster genom att kryssa för <span class="gui">Visa dolda filer</span>, från menyn <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="Visningsalternativ"></span></span> i verktygsfältet.</p>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div id="icon-view-defaults" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Standard för ikonvyn</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Förvald zoomnivå</span></dt>
<dd class="terms">
<p class="p">Du kan förstora eller förminska ikoner och text i ikonvyn med det här alternativet. Du kan också ändra den här inställningen i en individuell mapp genom att klicka på knappen <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="Visningsalternativ"></span></span> i verktygsfältet och välja <span class="gui">Zooma in</span>, <span class="gui">Zooma ut</span> eller <span class="gui">Normal storlek</span>. Om du ofta använder en större eller mindre zoomnivå kan du ange standarden med det här alternativet.</p>
<p class="p">I ikonvyn visas olika mängd <span class="link"><a href="nautilus-display.html#icon-captions" title="Ikontext">ikontext</a></span> baserat på din zoomnivå.</p>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div id="list-view-defaults" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Standard för listvy</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Förvald zoomnivå</span></dt>
<dd class="terms"><p class="p">Du kan förstora eller förminska ikoner och text i listvyn med det här alternativet. Du kan också ändra den här inställningen i en individuell mapp genom att klicka på knappen <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="Visningsalternativ"></span></span> i verktygsfältet och välja <span class="gui">Zooma in</span>, <span class="gui">Zooma ut</span> eller <span class="gui">Normal storlek</span>. Om du ofta använder en större eller mindre zoomnivå kan du ange standarden emd det här alternativet.</p></dd>
</dl></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="nautilus-prefs.html" title="Inställningar för filhanterare">Inställningar för filhanterare</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
