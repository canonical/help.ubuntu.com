<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Kolumninställningar för listvy i Filer</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 23.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a> » <a class="trail" href="nautilus-prefs.html.sv" title="Inställningar för filhanterare">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Kolumninställningar för listvy i Filer</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Det finns flera kolumner med information som du kan visa i listvyn i <span class="gui">Filer</span>. Högerklicka på en kolumnrubrik och markera eller avmarkera vilka kolumner som ska vara synliga.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Namn</span></dt>
<dd class="terms">
<p class="p">Namnet på mappar och filer.</p>
<div class="note note-tip" title="Tips">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m12 2c-3.8541 0-7 3.1459-7 7 0 1.823 0.4945 3.139 1.1641 4.133 0.6695 0.994 1.4328 1.671 2.039 2.471 0.0882 0.116 0.1749 0.656 0.2071 1.32 0.016 0.332 0.0133 0.68 0.1894 1.119 0.0881 0.22 0.2439 0.478 0.5059 0.672 0.2619 0.194 0.6028 0.285 0.8945 0.285h4c0.583 0 1.204-0.478 1.402-0.908 0.199-0.43 0.217-0.793 0.244-1.137 0.056-0.688 0.138-1.319 0.211-1.441 0.549-0.916 1.304-2.009 1.94-3.114 0.636-1.104 1.203-2.199 1.203-3.4 0-3.8541-3.146-7-7-7zm0 2c2.773 0 5 2.2267 5 5 0 0.456-0.359 1.401-0.936 2.402-0.111 0.195-0.246 0.399-0.369 0.598h-7.8825c-0.4871-0.728-0.8125-1.519-0.8125-3 0-2.7733 2.2267-5 5-5z" style="block-progression:tb;color-rendering:auto;color:#000000;image-rendering:auto;isolation:auto;mix-blend-mode:normal;shape-rendering:auto;solid-color:#000000;text-decoration-color:#000000;text-decoration-line:none;text-decoration-style:solid;text-indent:0;text-transform:none;white-space:normal"></path>
 <path class="yelp-svg-fill" d="m9 20a0.5 0.5 0 0 0-0.5 0.5 0.5 0.5 0 0 0 0.5 0.5h6a0.5 0.5 0 0 0 0.5-0.5 0.5 0.5 0 0 0-0.5-0.5h-6zm0 2a0.5 0.5 0 0 0-0.5 0.5 0.5 0.5 0 0 0 0.5 0.5h6a0.5 0.5 0 0 0 0.5-0.5 0.5 0.5 0 0 0-0.5-0.5h-6z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p"><span class="gui">Namn</span>-kolumnen kan inte gömmas.</p></div></div></div>
</div>
</dd>
<dt class="terms"><span class="gui">Storlek</span></dt>
<dd class="terms"><p class="p">Storleken för en mapp anges som antalet av objekt som finns i mappen. Storleken för en fil anges som byte, KB, eller MB.</p></dd>
<dt class="terms"><span class="gui">Typ</span></dt>
<dd class="terms"><p class="p">Visas som mapp, eller filtyp som PDF-dokument, JPEG-bild, MP3-ljud, med mera.</p></dd>
<dt class="terms"><span class="gui">Ändrad</span></dt>
<dd class="terms"><p class="p">Visar datum då filen senast ändrades.</p></dd>
<dt class="terms"><span class="gui">Ägare</span></dt>
<dd class="terms"><p class="p">Namnet på användaren som äger filen eller mappen.</p></dd>
<dt class="terms"><span class="gui">Grupp</span></dt>
<dd class="terms"><p class="p">Gruppen som äger filen. Varje användare är normalt i sin egen grupp, men det är möjligt att ha många användare i en grupp. En avdelning kan till exempel ha en egen grupp i en arbetsmiljö.</p></dd>
<dt class="terms"><span class="gui">Rättigheter</span></dt>
<dd class="terms">
<p class="p">Visar filrättigheterna. Till exempel <span class="gui">drwxrw-r--</span></p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Det första tecknet är filtypen. <span class="gui">-</span> innebär en normal fil och <span class="gui">d</span> innebär en mapp. I ovanliga fall kan andra tecken också visas.</p></li>
<li class="list"><p class="p">Nästa tre tecken <span class="gui">rwx</span> anger rättigheter för användaren som äger filen.</p></li>
<li class="list"><p class="p">Nästa tre <span class="gui">rw-</span> anger rättigheter för alla medlemmar i gruppen som äger filen.</p></li>
<li class="list"><p class="p">De sista tre tecknen i kolumnen <span class="gui">r--</span> ange rättigheter för alla andra användare på systemet.</p></li>
</ul></div></div></div>
<p class="p">Varje rättighet har följande innebörd:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p"><span class="gui">r</span>: läsbar, innebär att du kan öppna filen eller mappen</p></li>
<li class="list"><p class="p"><span class="gui">w</span>: skrivbar, innebär att du kan spara ändringar till den</p></li>
<li class="list"><p class="p"><span class="gui">x</span>: körbar, innebär att du kan köra den om det är program- eller skriptfil eller så kan du komma åt undermappar om det är en mapp</p></li>
<li class="list"><p class="p"><span class="gui">-</span>: rättighet inte inställd</p></li>
</ul></div></div></div>
</dd>
<dt class="terms"><span class="gui">MIME-typ</span></dt>
<dd class="terms"><p class="p">Visar objektets MIME-typ.</p></dd>
<dt class="terms"><span class="gui">Plats</span></dt>
<dd class="terms"><p class="p">Sökvägen till platsen för filen.</p></dd>
<dt class="terms"><span class="gui">Ändrad — Tid</span></dt>
<dd class="terms"><p class="p">Visar tid och datum då filen senast ändrades.</p></dd>
<dt class="terms"><span class="gui">Åtkommen</span></dt>
<dd class="terms"><p class="p">Visar tid eller datum då filen senast ändrades.</p></dd>
</dl></div></div></div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="nautilus-prefs.html.sv" title="Inställningar för filhanterare">Inställningar för filhanterare</a><span class="desc"> — Visa och ställ in inställningar för filhanteraren.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
