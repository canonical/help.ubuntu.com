<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Färghantering</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Färghantering</span></h1></div>
<div class="region">
<div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="color-assignprofiles.html.sv" title="Hur associerar jag färgprofiler till enheter?"><span class="title">Hur associerar jag färgprofiler till enheter?</span><span class="linkdiv-dash"> — </span><span class="desc">I <span class="guiseq"><span class="gui">Inställningar</span> ▸ <span class="gui">Färg</span></span> kan du lägga till en färgprofil för din skärm.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-whyimportant.html.sv" title="Varför är färghantering viktigt?"><span class="title">Varför är färghantering viktigt?</span><span class="linkdiv-dash"> — </span><span class="desc">Färghantering är viktigt för designers, fotografer och konstnärer.</span></a></div>
</div></div></div></div></div>
<section id="profiles"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Färgprofiler</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="color-howtoimport.html.sv" title="Hur importerar jag färgprofiler?"><span class="title">Hur importerar jag färgprofiler?</span><span class="linkdiv-dash"> — </span><span class="desc">Färgprofiler kan importeras genom att öppna dem.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-whatisprofile.html.sv" title="Vad är en färgprofil?"><span class="title">Vad är en färgprofil?</span><span class="linkdiv-dash"> — </span><span class="desc">En färgprofil är en enkel fil som visar en färgrymd eller hur en enhet svarar på färger.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="color-whatisspace.html.sv" title="Vad är en färgrymd?"><span class="title">Vad är en färgrymd?</span><span class="linkdiv-dash"> — </span><span class="desc">En färgrymd är ett definierat intervall av färger.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-gettingprofiles.html.sv" title="Var får jag tag på färgprofiler?"><span class="title">Var får jag tag på färgprofiler?</span><span class="linkdiv-dash"> — </span><span class="desc">Färgprofiler tillhandahålls av tillverkare men du kan också generera dem själv.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="calibration"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Kalibrering</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="color-calibrate-scanner.html.sv" title="Hur kalibrerar jag min bildläsare?"><span class="title">Hur kalibrerar jag min bildläsare?</span><span class="linkdiv-dash"> — </span><span class="desc">Att kalibrera din bildläsare är viktigt för att fånga korrekta färger.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-calibrate-camera.html.sv" title="Hur kalibrerar jag min kamera?"><span class="title">Hur kalibrerar jag min kamera?</span><span class="linkdiv-dash"> — </span><span class="desc">Att kalibrera din kamera är viktigt för att fånga korrekta färger.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-calibrate-printer.html.sv" title="Hur kalibrerar jag min skrivare?"><span class="title">Hur kalibrerar jag min skrivare?</span><span class="linkdiv-dash"> — </span><span class="desc">Det är viktigt att kalibrera din skrivare för att utskriften ska ge rätt färger.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-calibrate-screen.html.sv" title="Hur kalibrerar jag min skärm?"><span class="title">Hur kalibrerar jag min skärm?</span><span class="linkdiv-dash"> — </span><span class="desc">Att kalibrera din skärm är viktigt för att visa korrekta färger.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-canshareprofiles.html.sv" title="Kan jag dela min färgprofil?"><span class="title">Kan jag dela min färgprofil?</span><span class="linkdiv-dash"> — </span><span class="desc">Att dela färgprofiler är aldrig en bra idé eftersom hårdvara förändras över tid.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="color-calibrationcharacterization.html.sv" title="Vad är skillnaden mellan kalibrering och karakterisering?"><span class="title">Vad är skillnaden mellan kalibrering och karakterisering?</span><span class="linkdiv-dash"> — </span><span class="desc">Kalibrering och karakterisering är helt olika saker.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-why-calibrate.html.sv" title="Varför måste jag själv kalibrera?"><span class="title">Varför måste jag själv kalibrera?</span><span class="linkdiv-dash"> — </span><span class="desc">Kalibrering är viktigt om du bryr dig om färgerna du visar eller skriver ut.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-calibrationdevices.html.sv" title="Vilka färgmätningsinstrument finns det stöd för?"><span class="title">Vilka färgmätningsinstrument finns det stöd för?</span><span class="linkdiv-dash"> — </span><span class="desc">Vi har stöd för ett stort antal kalibreringsenheter.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-calibrationtargets.html.sv" title="Vilka måltyper finns det stöd för?"><span class="title">Vilka måltyper finns det stöd för?</span><span class="linkdiv-dash"> — </span><span class="desc">Kalibreringsmål behövs för att genomföra profilering av bildläsare och kamera.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="problems"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Problem</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="color-testing.html.sv" title="Hur testar jag om färghanteringen fungerar korrekt?"><span class="title">Hur testar jag om färghanteringen fungerar korrekt?</span><span class="linkdiv-dash"> — </span><span class="desc">Använd de tillhandahållna profilerna för att kontrollera att dina profiler appliceras korrekt för din skärm.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-notifications.html.sv" title="Kan jag bli aviserad när min färgprofil är felaktig?"><span class="title">Kan jag bli aviserad när min färgprofil är felaktig?</span><span class="linkdiv-dash"> — </span><span class="desc">Du kan bli aviserad om din färgprofil är gammal och otillförlitlig.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="color-missingvcgt.html.sv" title="Saknas information för helskärmsfärgkalibrering?"><span class="title">Saknas information för helskärmsfärgkalibrering?</span><span class="linkdiv-dash"> — </span><span class="desc">Helskärmsfärgkorrigering modifierar alla skärmfärger för alla fönster.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="color-notspecifiededid.html.sv" title="Varför har inte standardprofilerna för skärmar ett utgångsdatum?"><span class="title">Varför har inte standardprofilerna för skärmar ett utgångsdatum?</span><span class="linkdiv-dash"> — </span><span class="desc">Standardprofiler för skärmar har inget kalibreringsdatum.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — Få GNOME att arbeta för dig, från hårdvarukontroll till sekretessinställningar.</span>
</li>
<li class="links ">
<a href="hardware.html.sv" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a><span class="desc"> — Konfigurera hårdvara och diagnostisera problem, inklusive skrivare, skärmar, diskar med mera.</span>
</li>
</ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
