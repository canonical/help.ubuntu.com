<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Dokument</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#documents" title="Dokument">Dokument</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Dokument</span></h1></div>
<div class="region">
<div class="contents"><p class="p"><span class="app">Dokument</span> är ett GNOME-program som låter dig visa, organisera, och skriva ut dokument på din dator eller som skapats via internet med <span class="em">Google Docs</span> eller <span class="em">SkyDrive</span>.</p></div>
<div id="view" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Visa, sortera och sök</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="documents-formats.html" title="Format som stöds"><span class="title">Format som stöds</span><span class="linkdiv-dash"> — </span><span class="desc"><span class="app">Dokument</span> visar ett antal populära dokumenttyper.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="documents-view.html" title="Visa dokument som lagras lokalt eller online"><span class="title">Visa dokument som lagras lokalt eller online</span><span class="linkdiv-dash"> — </span><span class="desc">Visa dokument över hela skärmen.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="documents-filter.html" title="Filtrera dokument"><span class="title">Filtrera dokument</span><span class="linkdiv-dash"> — </span><span class="desc">Välj vilka dokument du vill visa.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="documents-search.html" title="Sök efter filer"><span class="title">Sök efter filer</span><span class="linkdiv-dash"> — </span><span class="desc">Hitta rätt dokument genom att leta efter titel eller författare.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="documents-viewgrid.html" title="Visa filer i en lista eller ett rutnät"><span class="title">Visa filer i en lista eller ett rutnät</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra hur dokument visas.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="documents-info.html" title="Hitta information om dokument"><span class="title">Hitta information om dokument</span><span class="linkdiv-dash"> — </span><span class="desc">Se ett dokuments namn, plats, ändringsdatum, eller typ.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="print" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Välj, sortera, skriv ut</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="documents-collections.html" title="Gör samlingar av dokument"><span class="title">Gör samlingar av dokument</span><span class="linkdiv-dash"> — </span><span class="desc">Gruppera relaterade dokument i en samling.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="documents-select.html" title="Markera dokument"><span class="title">Markera dokument</span><span class="linkdiv-dash"> — </span><span class="desc">Använd markeringsläget till att välja fler än ett dokument eller samling.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="documents-print.html" title="Skriv ut ett dokument"><span class="title">Skriv ut ett dokument</span><span class="linkdiv-dash"> — </span><span class="desc">Skriv ut dokument som lagras lokalt eller online.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="question" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Frågor</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="documents-tracker.html" title="Mina dokument syns inte"><span class="title">Mina dokument syns inte</span><span class="linkdiv-dash"> — </span><span class="desc">Lokala eller fjärrdokument visas inte.</span></a></div></div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="documents-previews.html" title="Varför har inte somliga filer någon förhandsgranskning?"><span class="title">Varför har inte somliga filer någon förhandsgranskning?</span><span class="linkdiv-dash"> — </span><span class="desc">Du kan bara förhandsgranska filer som lagras lokalt.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html#documents" title="Dokument">Dokument</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
