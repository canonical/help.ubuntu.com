<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Anslut din dator till en Bluetooth-enhet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="bluetooth.html" title="Bluetooth">Bluetooth</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Anslut din dator till en Bluetooth-enhet</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Innan du kan använda en Bluetooth-enhet, som en mus eller ett par hörlurar, måste du först ansluta din dator till enheten. Detta kallas också att para Bluetooth-enheterna.</p>
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">Innan du börjar, se till att Bluetooth är aktiverat på din dator. Se <span class="link"><a href="bluetooth-turn-on-off.html" title="Bluetooth på/av">Bluetooth på/av</a></span>.</p></div></div></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på Bluetooth-ikonen i menyraden och välj <span class="gui">Ställ in ny enhet</span>.</p></li>
<li class="steps"><p class="p">Gör den andra Bluetooth-enheten <span class="link"><a href="bluetooth-visibility.html" title="Vad är Bluetooth-synlighet?">upptäckbar, eller synlig</a></span>, och placera den inom 10 meters avstånd från din dator. Klicka på <span class="gui">Fortsätt</span>. Din dator kommer börja leta efter enheter.</p></li>
<li class="steps"><p class="p">Om för många enheter hittas, använd den utfällbara menyn <span class="gui">Enhetstyp</span> för att bara visa en viss typ av enhet i listan.</p></li>
<li class="steps">
<p class="p">Klicka på <span class="gui">PIN-alternativ</span> för att ange hur en PIN-kod ska levereras till den andra enheten.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Den automatiska PIN-inställningen kommer använda en sexsiffrig numerisk kod. En enhet utan tangenter eller skärm, som en mus eller ett headset, kan kräva en specifik PIN-kod, som 0000, eller ingen PIN-kod alls. Se enhetens manual för korrekt inställning.</p></div></div></div></div>
<p class="p">Välj en lämplig PIN-inställning för din enhet, och klicka sedan på <span class="gui">Stäng</span>.</p>
</li>
<li class="steps"><p class="p">Klicka på <span class="gui">Fortsätt</span> för att fortsätta. Om du inte valde ett förvalt PIN kommer PIN-koden visas på skärmen.</p></li>
<li class="steps">
<p class="p">Om det behövs, bekräfta PIN-koden på din andra enhet. Enheten bör visa dig PIN-koden du ser på din dators skärm, eller be dig mata in PIN-koden. Bekräfta PIN-koden på enheten och klicka sedan på <span class="gui">Stämmer</span>.</p>
<p class="p">Du måste slutföra inmatningen inom 20 sekunder på de flesta enheter, annars släpps anslutningen. Om det händer, gå tillbaka till enhetslistan och börja om från början.</p>
</li>
<li class="steps"><p class="p">Ett meddelande visas när anslutningen etableras. Klicka på <span class="gui">Stäng</span>.</p></li>
</ol></div></div></div>
<p class="p">Du kan <span class="link"><a href="bluetooth-remove-connection.html" title="Ta bort en anslutning mellan Bluetooth-enheter">ta bort en Bluetooth-anslutning</a></span> vid ett senare tillfälle, om så önskas.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">För att ha kontroll över åtkomst till dina delade filer, se inställningarna för <span class="gui">Bluetooth-delning</span>. Se <span class="link"><a href="sharing-bluetooth.html" title="Styr delning över Bluetooth">Styr delning över Bluetooth</a></span>.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="bluetooth.html" title="Bluetooth">Bluetooth</a><span class="desc"> — <span class="link"><a href="bluetooth-connect-device.html" title="Anslut din dator till en Bluetooth-enhet">Anslut</a></span>, <span class="link"><a href="bluetooth-send-file.html" title="Skicka en fil till en Bluetooth-enhet">skicka filer</a></span>, <span class="link"><a href="bluetooth-turn-on-off.html" title="Bluetooth på/av">slå på och av</a></span>...</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="sharing-bluetooth.html" title="Styr delning över Bluetooth">Styr delning över Bluetooth</a><span class="desc"> — Alternativ för Bluetooth-fildelning och -mottagande.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
