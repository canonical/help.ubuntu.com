<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Qemu</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="virtualization.html" title="Virtualisering">Virtualisering</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="libvirt.html" title="libvirt">Föregående</a><a class="nextlinks-next" href="cloud-images-and-uvtool.html" title="Cloud images and uvtool">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Qemu</h1></div>
<div class="region">
<div class="contents">
<p class="para">
        <a href="http://wiki.qemu.org/Main_Page" class="ulink" title="http://wiki.qemu.org/Main_Page">Qemu</a> is a machine emulator that can run operating systems and programs for one machine on a different machine.
        Mostly it is not used as emulator but as virtualizer in collaboration with KVM or XEN kernel components. In that case it utilizes the virtualization technology of the hardware to virtualize guests.
    </p>
<p class="para">
        While qemu has a <a href="http://wiki.qemu.org/download/qemu-doc.html#sec_005finvocation" class="ulink" title="http://wiki.qemu.org/download/qemu-doc.html#sec_005finvocation">command line interface</a> and a <a href="http://wiki.qemu.org/download/qemu-doc.html#pcsys_005fmonitor" class="ulink" title="http://wiki.qemu.org/download/qemu-doc.html#pcsys_005fmonitor">monitor</a> to interact with running guests those is rarely used that way for other means than development purposes.
        <a class="link" href="libvirt.html" title="libvirt">Libvirt</a> provides an abstraction from specific versions and hypervisors and encapsulates some workarounds and best practices.
    </p>
</div>
<div class="links sectionlinks" role="navigation"><ul><li class="links"><a class="xref" href="qemu.html#machine-type-upgrade" title="Upgrading the machine type">Upgrading the machine type</a></li></ul></div>
<div class="sect2 sect" id="machine-type-upgrade"><div class="inner">
<div class="hgroup"><h2 class="title">Upgrading the machine type</h2></div>
<div class="region"><div class="contents">
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="para">This also is documented along some more constraints and considerations at the <a href="https://wiki.ubuntu.com/QemuKVMMigration#Upgrade_machine_type" class="ulink" title="https://wiki.ubuntu.com/QemuKVMMigration#Upgrade_machine_type">Ubuntu Wiki</a></p></div></div></div></div>
<p class="para">You might want to update your machine type of an existing defined guest to:</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist"><p class="para">to pick up latest security fixes and features</p></li>
<li class="list itemizedlist"><p class="para">continue using a guest created on a now unsupported release</p></li>
</ul></div>
<p class="para">In general it is recommended to update machine types when upgrading qemu/kvm to a new major version. But this can likely never be an automated task as this change is guest visible. The guest devices might change in appearance, new features will be announced to the guest and so on. Linux is usually very good at tolerating such changes, but it depends so much on the setup and workload of the guest that this has to be evaluated by the owner/admin of the system. Other operating systems where known to often have severe impacts by changing the hardware. Consider a machine type change similar to replacing all devices and firmware of a physical machine to the latest revision - all considerations that apply there apply to evaluating a machine type upgrade as well.</p>
<p class="para">As usual with major configuration changes it is wise to back up your guest definition and disk state to be able to do a rollback just in case. There is no integrated single command to update the machine type via virsh or similar tools. It is a normal part of your machine definition. And therefore updated the same way as most others.</p>
<p class="para">First shutdown your machine and wait until it has reached that state.</p>
<div class="screen"><pre class="contents ">virsh shutdown &lt;yourmachine&gt;
# wait
virsh list --inactive
# should now list your machine as "shut off"
        </pre></div>
<p class="para">Then edit the machine definition and find the type in the type tag at the machine attribute.</p>
<div class="screen"><pre class="contents ">virsh edit &lt;yourmachine&gt;
&lt;type arch='x86_64' machine='pc-i440fx-xenial'&gt;hvm&lt;/type&gt;
        </pre></div>
<p class="para">Change this to the value you want. If you need to check what types are available via "-M ?" Note that while providing upstream types as convenience only Ubuntu types are supported. There you can also see what the current default would be. In general it is strongly recommended that you change to newer types if possible to exploit newer features, but also to benefit of bugfixes that only apply to the newer device virtualization.</p>
<div class="screen"><pre class="contents ">kvm -M ?
# lists machine types, e.g.
pc-i440fx-xenial       Ubuntu 16.04 PC (i440FX + PIIX, 1996) (default)
...
        </pre></div>
<p class="para">After this you can start your guest again. You can check the current machine type from guest and host depending on your needs.</p>
<div class="screen"><pre class="contents ">virsh start &lt;yourmachine&gt;
# check from host, via dumping the active xml definition
virsh dumpxml &lt;yourmachine&gt; | xmllint --xpath "string(//domain/os/type/@machine)" -
# or from the guest via dmidecode
sudo dmidecode | grep Product -A 1
        Product Name: Standard PC (i440FX + PIIX, 1996)
        Version: pc-i440fx-xenial
        </pre></div>
<p class="para">If you keep non-live definitions around like xml files remember to update those as well.</p>
</div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="libvirt.html" title="libvirt">Föregående</a><a class="nextlinks-next" href="cloud-images-and-uvtool.html" title="Cloud images and uvtool">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
