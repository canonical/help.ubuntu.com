<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skriva ut kuvert</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="printing.html" title="Utskrifter">Utskrifter</a> › <a class="trail" href="printing.html#paper" title="Olika pappersstorlekar och layouter">Storlekar och layouter</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Skriva ut kuvert</span></h1></div>
<div class="region">
<div class="contents"><p class="p">De flesta skrivare låter dig skriva ut direkt på ett kuvert. Detta är särskilt användbart om du till exempel har många brev att skicka.</p></div>
<div id="envelope" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Skriva ut på kuvert</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Det finns två saker du måste kontrollera när du försöker att skriva ut på ett kuvert.</p>
<p class="p">Det första är att din skrivare vet vilken storlek kuvertet har. Tryck på <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>P</kbd></span></span> för att öppna utskriftsdialogen, gå till fliken <span class="gui">Sidinställning</span> och som <span class="gui">Papperstyp</span> välj ”Kuvert” om du kan. Om du inte kan göra detta, se om du kan ändra <span class="gui">Pappersstorlek</span> till en kuvertstorlek (till exempel <span class="gui">C5</span>). På bunten med kuvert bör det stå vilken storlek de har; de flesta kuvert levereras i standardstorlekar.</p>
<p class="p">För det andra måste du säkerställa att kuverten matas in med rätt sida upp i skrivaren. Kontrollera skrivarens manual för hur du gör detta eller försök att skriva ut ett enstaka kuvert och kontrollera vilken sida som skrivs ut på för att se vilket håll som ska vara uppåt.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">Vissa skrivare är inte designade för att kunna skriva ut kuvert, speciellt vissa laserskrivare. Kontrollera din skrivares manual för att se om den kan skriva ut på kuvert. Annars kan du skada skrivaren genom att mata in ett kuvert.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="printing.html#paper" title="Olika pappersstorlekar och layouter">Olika pappersstorlekar och layouter</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
