<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Fönsteråtgärder</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord</a> › <a class="trail" href="shell-overview.html#apps" title="Program och fönster">Program och fönster</a> » <a class="trail" href="shell-windows.html" title="Fönster och arbetsytor">Fönster och arbetsytor</a> › <a class="trail" href="shell-windows.html#working-with-windows" title="Arbeta med fönster">Fönster</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Fönsteråtgärder</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Du kan ändra storlek på eller gömma fönster för att bättre passa ditt arbetsflöde.</p></div>
<div id="min-rest-close" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Minimera, återställ och stäng</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att minimera eller dölja ett fönster:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">Klicka på <span class="gui">-</span> längst upp till vänster i programmets <span class="gui">menyrad</span>. Om programmet är maximerat (tar upp hela skärmen) kommer menyraden visas längst upp i skärmen. Annars finns minimeraknappen längst upp i programmets fönster.</p></li>
<li class="list"><p class="p">Eller tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span> för att öppna fönstermenyn. Tryck sedan <span class="key"><kbd>n</kbd></span>. Fönstret "försvinner" in i Startaren.</p></li>
</ul></div></div></div>
<p class="p">För att återställa fönstret:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc"><li class="list"><p class="p">Klicka på det i <span class="link"><a href="unity-launcher-intro.html" title="Använda programstartaren">Startaren</a></span> eller leta fram det i fönsterväxlaren genom att trycka <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span>.</p></li></ul></div></div></div>
<p class="p">För att stänga fönstret:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">Klicka på <span class="gui">x</span>:et längst upp till vänster i fönstret, eller</p></li>
<li class="list"><p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F4</kbd></span></span> eller</p></li>
<li class="list"><p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span> för att öppna fönstermenyn. Tryck sedan <span class="key"><kbd>t</kbd></span>.</p></li>
</ul></div></div></div>
</div></div>
</div></div>
<div id="resize" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ändra storlek</span></h2></div>
<div class="region"><div class="contents">
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan inte ändra ett fönsters storlek om det är <span class="em">maximerat</span>.</p></div></div></div></div>
<p class="p">För att ändra fönsterstorlek horisontellt och/eller vertikalt:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc"><li class="list"><p class="p">Flytta muspekaren till något av fönstrets hörn tills den ändras till en "hörnpekare". Klicka, håll, och dra för att ändra fönsterstorleken i valfri riktning.</p></li></ul></div></div></div>
<p class="p">För att bara ändra horisontell storlek:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc"><li class="list"><p class="p">Flytta muspekaren till endera sida av fönstret tills den ändras till en "sidopekare". Klicka, håll, och dra för att ändra fönstrets horisontella storlek.</p></li></ul></div></div></div>
<p class="p">För att bara ändra vertikal storlek:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc"><li class="list"><p class="p">Flytta muspekaren till fönstrets topp eller bas tills den ändras till en "toppekare" respektive "bottenpekare". Klicka, håll, och dra för att ändra fönstrets vertikala storlek.</p></li></ul></div></div></div>
</div></div>
</div></div>
<div id="arrange" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ordna fönster på din arbetsyta</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att placera två fönster bredvid varandra:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ett fönsters <span class="gui">titellist</span> och dra den mot skärmens vänstra kant. När <span class="gui">muspekaren</span> når kanten kommer skärmens vänstra halva markeras. Släpp musknappen, så kommer fönstret fylla skärmens vänstra halva.</p></li>
<li class="steps"><p class="p">Dra ett annat fönster till höger: när skärmens högra halva är markerad, släpp. De båda fönstren fyller nu varsin halva av skärmen.</p></li>
</ol></div></div></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du trycker <span class="key"><kbd>Alt</kbd></span> och sedan klickar varsomhelst i ett fönster kan du flytta fönstret. Vissa upplever det här som lättare än att klicka på ett programs <span class="gui">titellist</span>.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-windows.html#working-with-windows" title="Arbeta med fönster">Arbeta med fönster</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links "><a href="unity-menubar-intro.html#window-management" title="Fönsterhanteringsknappar">Fönsterhanteringsknappar</a></li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
