<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Öppna filer med andra program</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Öppna filer med andra program</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">När du dubbelklickar på en fil i filhanteraren kommer den öppnas med det förvalda programmet för den filtypen. Du kan öppna den i ett annat program, söka på internet efter program, eller ange ett förvalt program för alla filer av den typen.</p>
<p class="p">För att öppna en fil med ett program annat än det förvalda, högerklicka på filen och välj programmet du vill starta från menyns övre del. Om du inte ser programmet du vill ha, klicka på <span class="gui">Öppna med annat program</span>. Som standard visar filhanteraren bara program som den vet kan arbeta med filen. För att gå igenom alla program på din dator, klicka på <span class="gui">Visa andra program</span>.</p>
<p class="p">Om du fortfarande inte kan hitta rätt program kan du söka efter fler program genom att klicka på <span class="gui">Hitta program på nätet</span>. Filhanteraren kommer då söka på internet efter paket som innehåller program som man vet kan arbeta med filer av den typen.</p>
</div>
<div id="default" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ändra förvalt program</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan ändra vilket program som ska vara förvalt när filer av en viss typ öppnas. Detta låter dig öppna ditt favoritprogram när du dubbelklickar för att öppna en fil. Du kan till exempel vilja att din favoritmusikspelare öppnas när du dubbelklickar på en MP3-fil.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Välj en fil av den typ vars förvalda program du vill ändra. För att ändra vilket program används för att öppna till exempel MP3-filer, välj en <span class="file">.mp3</span>-fil.</p></li>
<li class="steps"><p class="p">Högerklicka på filen och välj <span class="gui">Egenskaper</span>.</p></li>
<li class="steps"><p class="p">Välj fliken <span class="gui">Öppna med</span>.</p></li>
<li class="steps">
<p class="p">Välj programmet du önskar och klicka <span class="gui">Ange som standard</span>. Som standard visar filhanteraren endast program som den vet kan hantera filen. För att leta genom alla program på din dator, klicka på <span class="gui">Visa andra program</span>.</p>
<p class="p">Om <span class="gui">Andra program</span> innehåller ett program som du ibland vill använda, men inte som förval, välj programmet och klicka på <span class="gui">Lägg till</span>. Detta lägger till programmet i <span class="gui">Rekommenderade program</span>. Du kommer sedan kunna använda det här programmet genom att högerklicka på filen och välja det från listan.</p>
</li>
</ol></div></div></div>
<p class="p">Detta ändrar förvalt program inte bara för den valda filen, utan för alla filer av samma typ.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
