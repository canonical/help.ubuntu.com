<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Filhanterarens visningsinställningar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#more-file-tasks" title="Fler filrelaterade uppgifter">Fler filrelaterade uppgifter</a> » <a class="trail" href="nautilus-prefs.html" title="Inställningar för filhanterare">Inställningar för filhanterare</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Filhanterarens visningsinställningar</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Du kan styra hur filhanteraren visar text under ikoner. Klicka på <span class="gui">Filer</span> i systemraden, välj <span class="gui">Inställningar</span> och välj fliken <span class="gui">Visa</span>.</p></div>
<div id="icon-captions" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ikonrubriker</span></h2></div>
<div class="region"><div class="contents">
<div class="media media-image floatend"><div class="inner"><img src="figures/nautilus-icons.png" height="110" width="250" class="media media-block" alt="Filhanterarens ikoner med text"></div></div>
<p class="p">När du använder ikonvyn kan du välja att visa extra information om filer och mappar som en text under varje ikon. Detta är till exempel användbart om du ofta behöver se vem som äger en fil eller när den senast modifierades.</p>
<p class="p">Du kan zooma i en mapp genom att klicka på knappen visningsalternativ i verktygsfältet och välja en zoomnivå med skjutreglaget. När du zoomar in kommer filhanteraren att visa mer och mer information i rubriker. Du kan välja upp till tre saker att visa i rubrikerna. Den första kommer att visas på de flesta zoomnivåerna. Den sista kommer bara att visas vid väldigt stora storlekar.</p>
<p class="p">Informationen du kan visa i ikonrubriker är samma som kolumnerna du kan använda i listvyn. Se <span class="link"><a href="nautilus-list.html" title="Kolumninställningar för listvy i Filer">Kolumninställningar för listvy i Filer</a></span> för mer information.</p>
</div></div>
</div></div>
<div id="list-view" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Listvy</span></h2></div>
<div class="region"><div class="contents"><p class="p">När du tittar på filer som en lista kan du <span class="gui">Navigera mappar i ett träd</span>. Detta visar expanderare för varje katalog i fillistan så att innehållet för flera kataloger kan visas samtidigt. Detta är användbart om mappstrukturen är relevant, t.ex. om dina musikfiler är organiserade med en mapp per artist och en undermapp per album.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="nautilus-prefs.html" title="Inställningar för filhanterare">Inställningar för filhanterare</a><span class="desc"> — Visa och ställ in inställningar för filhanteraren.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
