<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Svara på meddelande</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Svara på meddelande</span></h1></div>
<div class="region">
<div class="contents"><div class="ui-tile ">
<a href="figures/gnome-responding-to-messages.webm" class="ui-overlay"><span class="ui-tile-img" style="width: 812px; height: 452px;"><img src="gs-thumb-responding-to-messages.svg" width="812" height="452"></span></a><div class="ui-overlay"><div class="inner">
<a href="#" class="ui-overlay-close" title="Stäng">⨯</a><div class="contents"><div class="media media-video"><div class="inner">
<video src="figures/gnome-responding-to-messages.webm" preload="auto" controls="controls" class="media media-block" height="394" width="700" data-play-label="Spela upp" data-pause-label="Paus"></video><div class="media-ttml">
<div class="media-ttml-node media-ttml-div" data-ttml-begin="1" data-ttml-end="3"><div class="media-ttml-node media-ttml-p" data-ttml-begin="1" data-ttml-end="3">Svarar på meddelande</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="3" data-ttml-end="6"><div class="media-ttml-node media-ttml-p" data-ttml-begin="3" data-ttml-end="6">Flytta din mus över chattmeddelandet som visas nära toppen på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="6" data-ttml-end="9"><div class="media-ttml-node media-ttml-p" data-ttml-begin="6" data-ttml-end="9">Börja skriva ditt svar. När du är klar, tryck på <span class="key"><kbd>Retur</kbd></span> och skicka svaret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="9" data-ttml-end="10"><div class="media-ttml-node media-ttml-p" data-ttml-begin="9" data-ttml-end="10">Stäng chattmeddelandet.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="12" data-ttml-end="14"><div class="media-ttml-node media-ttml-p" data-ttml-begin="12" data-ttml-end="14">Fördröjt svar</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="16" data-ttml-end="22"><div class="media-ttml-node media-ttml-p" data-ttml-begin="16" data-ttml-end="22">Ett chattmeddelande nära toppen av skärmen försvinner efter en stund om du inte flyttar din mus över meddelandet.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="22" data-ttml-end="24"><div class="media-ttml-node media-ttml-p" data-ttml-begin="22" data-ttml-end="24">För att få tillbaka ditt obesvarade meddelande, klicka på klockan i systemraden.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="24" data-ttml-end="26"><div class="media-ttml-node media-ttml-p" data-ttml-begin="24" data-ttml-end="26">Från aviseringslistan, välj ditt meddelande.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="26" data-ttml-end="28"><div class="media-ttml-node media-ttml-p" data-ttml-begin="26" data-ttml-end="28">Börja skriva ditt svar.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="32" data-ttml-end="35"><div class="media-ttml-node media-ttml-p" data-ttml-begin="32" data-ttml-end="35">För att visa aviseringslistan, tryck <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>+<span class="key"><kbd>V</kbd></span></span>
</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="35" data-ttml-end="41"><div class="media-ttml-node media-ttml-p" data-ttml-begin="35" data-ttml-end="41">Använd piltangenterna för att välja meddelandet som du vill svara på, och tryck på <span class="key"><kbd>Retur</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="41" data-ttml-end="44"><div class="media-ttml-node media-ttml-p" data-ttml-begin="41" data-ttml-end="44">Börja skriva ditt svar.</div></div>
</div>
</div></div></div>
</div></div>
</div></div>
<div id="respond-to-messages-mouse" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Svara på ett chattmeddelande med musen</span></h2></div>
<div class="region"><div class="contents">
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Flytta din mus över chattmeddelandet som visas nära toppen på skärmen.</p></li>
<li class="steps"><p class="p">Börja skriv ditt svar och när du är klar, tryck på <span class="key"><kbd>Retur</kbd></span> för att skicka svaret.</p></li>
<li class="steps"><p class="p">För att stänga chattmeddelandet, klicka på stängknappen i det övre högra hörnet på chattmeddelandet.</p></li>
</ol></div></div></div>
<p class="p"></p>
</div></div>
</div></div>
<div id="respond-to-messages-delayed-mouse" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Fördröjt svar på ett chattmeddelande genom att använda musen</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">När ett chattmeddelande visas nära toppen på skärmen och du inte flyttar musen över meddelandet så kommer det att försvinna efter en stund.</p></li>
<li class="steps"><p class="p">För att få tillbaka ditt obesvarade meddelande, klicka på klockan i systemraden.</p></li>
<li class="steps"><p class="p">Från aviseringslistan, välj meddelandet du vill svara på och klicka på det.</p></li>
<li class="steps"><p class="p">När chattmeddelandet visas, börja skriva ditt svar.</p></li>
</ol></div></div></div></div></div>
</div></div>
<div id="respond-to-messages-delayed-keyboard" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Fördröjt svar på ett chattmeddelande genom att använda tangentbordet</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">För att få tillbaka ditt obesvarade chattmeddelande, tryck <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>+<span class="key"><kbd>V</kbd></span></span> för att visa listan över obesvarade aviseringar.</p></li>
<li class="steps"><p class="p">Använd piltangenterna för att välja aviseringen som du vill svara på, och tryck på <span class="key"><kbd>Retur</kbd></span>.</p></li>
<li class="steps"><p class="p">När chattmeddelandet visas, börja skriva ditt svar.</p></li>
</ol></div></div></div></div></div>
</div></div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p>You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
