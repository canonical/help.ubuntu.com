<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Välj ditt lösenord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="user-accounts.html" title="Användarkonton">Users</a> › <a class="trail" href="user-accounts.html#passwords" title="Lösenord">Lösenord</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Välj ditt lösenord</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">It is a good idea to change your password from time to time, especially if
  you think someone else knows what your password is.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Click the icon at the far right of the <span class="gui">menu bar</span> and select <span class="gui">System Settings</span>.</p></li>
<li class="steps"><p class="p">Open <span class="gui">User Accounts</span>.</p></li>
<li class="steps">
<p class="p">Click the label next to <span class="gui">Password</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">The label should look
    like a series of dots or boxes if you already have a password set.</p></div></div></div></div>
</li>
<li class="steps">
<p class="p">Enter your current password, then a new password. Enter your new
    password again in the <span class="gui">Confirm password</span> field.</p>
<p class="p">You can also click the button next to the
    <span class="gui">New password</span> field to select a randomly generated secure password.
    These passwords are hard for others to guess, but they can be hard to
    remember, so be careful.</p>
</li>
<li class="steps"><p class="p">Click <span class="gui">Change</span>.</p></li>
</ol></div></div></div>
<p class="p">Make sure you <span class="link"><a href="user-goodpassword.html" title="Välj ett säkert lösenord">choose a good password</a></span>.
  This will help to keep your user account safe.</p>
</div>
<div id="changepass" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Change the keyring password</span></h2></div>
<div class="region"><div class="contents">
<p class="p">If you change your login password, it may become out of sync with the
  <span class="em">keyring password</span>. The keyring keeps you from having to remember lots
  of different passwords by just requiring one <span class="em">master</span> password to access
  them all. If you change your user password (see above), your keyring password
  will remain the same as your old password.  To change the keyring
  password (to match your login password):</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Open the <span class="app">Passwords and Keys</span> application from
    the <span class="gui">Dash</span>.</p></li>
<li class="steps"><p class="p">In the <span class="gui">View</span> menu, ensure <span class="gui">By keyring</span> is
     checked.</p></li>
<li class="steps"><p class="p">In the sidebar under <span class="gui">Passwords</span>, right-click on
     <span class="gui">Login keyring</span> and select <span class="gui">Change Password</span>.</p></li>
<li class="steps"><p class="p">Enter your <span class="gui">Old Password</span>, followed by your new
     <span class="gui">Password</span>, and <span class="gui">Confirm</span> your new password by entering
     it again.</p></li>
<li class="steps"><p class="p">Click <span class="gui">OK</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="user-accounts.html#passwords" title="Lösenord">Lösenord</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="user-goodpassword.html" title="Välj ett säkert lösenord">Välj ett säkert lösenord</a><span class="desc"> — 
      Use longer, more complicated passwords.
    </span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
