<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vad är HUD?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord</a> › <a class="trail" href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Vad är HUD?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p"><span class="gui">HUD</span>, eller <span class="gui">Heads Up Display</span>, är ett sökbaserat alternativ till traditionella menyer och introducerades i Ubuntu 12.04 LTS.</p>
<p class="p">Vissa program, som <span class="link"><a href="https://apps.ubuntu.com/cat/applications/gimp" title="https://apps.ubuntu.com/cat/applications/gimp">Gimp</a></span> eller <span class="link"><a href="https://apps.ubuntu.com/cat/applications/inkscape" title="https://apps.ubuntu.com/cat/applications/inkscape">Inkscape</a></span>, har hundratals menyobjekt. Om du använder liknande program kanske du kommer ihåg namnet på ett menyobjekt, men inte hur du hittar det i menyerna.</p>
<p class="p">Att använda en sökruta kan vara mycket snabbare än att navigera igenom invecklade menyhierarkier. HUD kan också vara lättare att använda än vanliga menyer eftersom vissa kan ha svårigheter med att styra en muspekare med tillräcklig precision.</p>
</div>
<div id="use-the-hud" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Att använda HUD</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att testa HUD:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Tryck på <span class="key"><kbd>Alt</kbd></span> för att öppna HUD.</p></li>
<li class="steps"><p class="p">Börja skriva.</p></li>
<li class="steps"><p class="p">När du ser ett resultat som du vill köra, använd upp- och nertangenterna för att markera resultatet, och tryck sedan <span class="key"><kbd>Retur</kbd></span>, eller klicka på ditt önskade sökresultat.</p></li>
<li class="steps"><p class="p">Om du ändrar dig och vill lämna HUD, tryck <span class="key"><kbd>Alt</kbd></span> igen eller <span class="key"><kbd>Esc</kbd></span>. Du kan också klicka varsomhelst utanför HUD för att stänga den.</p></li>
</ol></div></div></div>
<p class="p">HUD håller reda på din sökhistorik, och justerar sökresultaten för att vara än mer behjälplig ju mer du använder den.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
