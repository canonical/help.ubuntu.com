<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använd gester på styrplattor och pekskärmar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 25.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 25.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Använd gester på styrplattor och pekskärmar</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Flerfingersgester kan användas på styrplattor och pekskärmar för systemnavigering, såväl som i program.</p>
<p class="p">Ett antal program kan använda gester. I <span class="app">Dokumentvisare</span> kan dokument zoomas och svepas undan med gester, och <span class="app">Bildvisare</span> låter dig zooma, rotera och panorera.</p>
</div>
<section id="system"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Systemomfattande gester</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="table"><div class="inner"><div class="region"><table class="table" style="border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-overview.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td>
<p class="p"><span class="em">Öppna översiktsvyn Aktiviteter och programvyn</span></p>
<p class="p">Placera tre fingrar på styrplattan eller pekskärmen och gör en gest uppåt för att öppna översiktsvyn Aktiviteter.</p>
<p class="p">För att öppna programvyn, placera tre fingrar och gör en gest uppåt igen.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-workspaces.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p"><span class="em">Växla arbetsyta</span></p>
<p class="p">Placera tre fingrar på styrplattan eller pekskärmen och gör en gest åt vänster eller höger.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-unfullscreen.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p"><span class="em">Lämna helskärmsläge</span></p>
<p class="p">På en pekskärm, dra neråt från den övre kanten för att lämna helskärmsläget för alla fönster.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-osk.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p"><span class="em">Ta fram skärmtangentbordet</span></p>
<p class="p">På en pekskärm, dra uppåt från den nedre kanten för att få upp <span class="link"><a href="keyboard-osk.html.sv" title="Använd ett skärmtangentbord">skärmtangentbordet</a></span>, om skärmtangentbordet är aktiverat.</p>
</td>
</tr>
</table></div></div></div></div></div>
</div></section><section id="apps"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Programgester</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="table"><div class="inner"><div class="region"><table class="table" style="border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-tap.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td>
<p class="p"><span class="em">Öppna ett objekt, starta ett program, spela en sång</span></p>
<p class="p">Tryck på ett objekt.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-hold.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p"><span class="em">Välj ett objekt och liståtgärder som kan utföras</span></p>
<p class="p">Tryck och håll under en eller två sekunder.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-scroll.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p"><span class="em">Rulla ytan på skärmen</span></p>
<p class="p">Dra: svep med ett finger som rör ytan.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-pinch-to-zoom.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p"><span class="em">Ändra zoomnivå för en vy (<span class="app">Kartor</span>, <span class="app">Foton</span>)</span></p>
<p class="p">Tvåfingernypning eller utsträckning: Rör vid ytan med två fingrar medan du rör dem närmre mot eller längre ifrån varandra.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="media"><span class="media media-image"><img src="figures/touch-rotate.svg" width="128" class="media media-inline" alt=""></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p"><span class="em">Rotera ett foto</span></p>
<p class="p">Tvåfingersrotation: Rör vid ytan med två fingrar och rotera.</p>
</td>
</tr>
</table></div></div></div></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus, styrplatta &amp; pekskärm</a><span class="desc"> — Justera beteendet hos pekdon så att de uppfyller dina personliga krav.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
