<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Klicka, dra eller rulla med styrplattan</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="mouse.html" title="Mus">Mus</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Klicka, dra eller rulla med styrplattan</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Du kan klicka, dubbelklicka, dra, och rulla med din styrplatta, utan att behöva separata fysiska knappar.</p></div>
<div id="clickordrag" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Klicka eller dra</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan klicka eller dra med hjälp av din styrplatta.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="em">Systemmenyn</span> <span class="media"><span class="media media-image"><img src="figures/system-devices-panel.svg" class="media media-inline" alt="Kugghjulsikon"></span></span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Öppna <span class="gui">Mus &amp; styrplatta</span>.</p></li>
<li class="steps"><p class="p">I avsnittet <span class="gui">Styrplatta</span>, markera <span class="gui">Tryck för att klicka</span>.</p></li>
</ol></div></div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">För att klicka, tryck lätt en gång (men inte i det nedre eller övre högra hörnet).</p></li>
<li class="list"><p class="p">För att dubbelklicka, tryck två gånger.</p></li>
<li class="list"><p class="p">För att dra ett objekt, dubbeltryck; men lyft inte fingret efteråt. Dra objektet dit du vill ha det, och lyft sedan fingret för att släppa.</p></li>
<li class="list"><p class="p">För att högerklicka, peka en gång i nedre högra hörnet.</p></li>
<li class="list"><p class="p">För att mittenklicka, peka en gång i övre högra hörnet.</p></li>
</ul></div></div></div>
</div></div>
</div></div>
<div id="twofingerscroll" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Tvåfingersrullning</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan rulla via din styrplatta genom att använda två fingrar.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="em">Systemmenyn</span> <span class="media"><span class="media media-image"><img src="figures/system-devices-panel.svg" class="media media-inline" alt="Kugghjulsikon"></span></span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Öppna <span class="gui">Mus &amp; styrplatta</span>.</p></li>
<li class="steps"><p class="p">I avsnittet <span class="gui">Styrplatta</span>, markera <span class="gui">Tvåfingersrullning</span>.</p></li>
</ol></div></div></div>
<p class="p">När det här väljs kommer trycka och dra med ett finger fungera som vanligt, men om du drar två fingrar över någon del av styrplattan kommer den rulla istället. Om du också väljer <span class="gui">Aktivera horisontell rullning</span> kan du röra dina fingrar till vänster och höger för att rulla horisontellt. Var noga med att hålla dina fingrar en bit isär. Om dina fingrar är för tätt ihop kan styrplattan känna av dem som ett enda stort finger.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Tvåfingersrullning kanske inte fungerar på alla styrplattor.</p></div></div></div></div>
</div></div>
</div></div>
<div id="contentsticks" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Innehåll fastnar vid fingrarna</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan dra innehåll som om du flyttade en fysisk bit papper via styrplattan.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="em">Systemmenyn</span> <span class="media"><span class="media media-image"><img src="figures/system-devices-panel.svg" class="media media-inline" alt="Kugghjulsikon"></span></span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Öppna <span class="gui">Mus &amp; styrplatta</span>.</p></li>
<li class="steps"><p class="p">I avsnittet <span class="gui">Styrplatta</span>, kryssa för <span class="gui">Innehåll fastnar vid fingrarna</span>.</p></li>
</ol></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Funktionen kallas också <span class="em">Naturlig rullning</span> eller <span class="em">Omvänd rullning</span>.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="mouse.html" title="Mus">Mus</a><span class="desc"> — <span class="link"><a href="mouse-lefthanded.html" title="Använd din mus med vänster hand">Vänsterhänt</a></span>, <span class="link"><a href="mouse-sensitivity.html" title="Justera hastigheten för musen och styrplattan">hastighet och känslighet</a></span>, <span class="link"><a href="mouse-touchpad-click.html" title="Klicka, dra eller rulla med styrplattan">styrplatteklick och rullning</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="unity-scrollbars-intro.html" title="Vad är överlagda rullningslister?">Vad är överlagda rullningslister?</a><span class="desc"> — Överlagda rullningslister är de tunna orange remsorna på långa dokument.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
