<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Inställningar för filhanterarens listkolumner</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » <a class="trail" href="nautilus-prefs.html" title="Inställningar för filhanterare">Inställningar för filhanterare</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Inställningar för filhanterarens listkolumner</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Det finns nio informationskolumner som du kan visa i filhanterarens listvy. Klicka på <span class="gui">Filer</span> i menyraden, välj <span class="gui">Inställningar</span> och välj fliken <span class="gui">Listkolumner</span> för att välja vilka kolumner som ska vara synliga.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Använd knapparna <span class="gui">Flytta upp</span> och <span class="gui">Flytta ner</span> för att bestämma i vilken ordning de markerade kolumnerna ska visas.</p></div></div></div></div>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Namn</span></dt>
<dd class="terms"><p class="p">Namnen på mappar och filer i den visade mappen.</p></dd>
<dt class="terms"><span class="gui">Storlek</span></dt>
<dd class="terms"><p class="p">Storleken på en mapp anges som antal objekt som finns i mappen. Filstorlek anges som byte, KB, eller MB.</p></dd>
<dt class="terms"><span class="gui">Typ</span></dt>
<dd class="terms"><p class="p">Visas som mapp, eller filtyp som PDF-dokument, JPEG-bild, MP3-ljud, med mera.</p></dd>
<dt class="terms"><span class="gui">Ändrad</span></dt>
<dd class="terms"><p class="p">Visar när filen senast ändrades.</p></dd>
<dt class="terms"><span class="gui">Ägare</span></dt>
<dd class="terms"><p class="p">Namn på användaren som äger mappen eller filen.</p></dd>
<dt class="terms"><span class="gui">Grupp</span></dt>
<dd class="terms"><p class="p">Gruppen som äger filen. På mina hemdatorer tillhör varje användare sin egen grupp. Grupper används ibland i företagsmiljöer, där användare kan sorteras in i grupper beroende på avdelningar eller projekt.</p></dd>
<dt class="terms"><span class="gui">Rättigheter</span></dt>
<dd class="terms">
<p class="p">Visar filåtkomsträttigheter, t.ex. <span class="gui">drwxrw-r--</span></p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">Det första tecknet, <span class="gui">d</span>, är filtypen. <span class="gui">-</span> betyder att det är en vanlig fil, och <span class="gui">d</span>betyder katalog (mapp).</p></li>
<li class="list"><p class="p">De tre följande tecknen <span class="gui">rwx</span> anger rättigheter för användaren som äger filen.</p></li>
<li class="list"><p class="p">Nästa tre <span class="gui">rw-</span> anger rättigheter för alla medlemmar i gruppen som äger filen.</p></li>
<li class="list"><p class="p">De sista tre tecknen i kolumnen <span class="gui">r--</span> anger rättigheter för alla andra användare på systemet.</p></li>
</ul></div></div></div>
<p class="p">Varje tecken har följande betydelser:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">r : Läsrättighet.</p></li>
<li class="list"><p class="p">w : Skrivrättighet.</p></li>
<li class="list"><p class="p">x : Körrättighet.</p></li>
<li class="list"><p class="p">- : Inga rättigheter.</p></li>
</ul></div></div></div>
</dd>
<dt class="terms"><span class="gui">MIME-typ</span></dt>
<dd class="terms"><p class="p">Visar objektets MIME-typ.</p></dd>
<dt class="terms"><span class="gui">Plats</span></dt>
<dd class="terms"><p class="p">Sökvägen till filens plats.</p></dd>
</dl></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="nautilus-prefs.html" title="Inställningar för filhanterare">Inställningar för filhanterare</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
