<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Installera från CD</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="installation.html" title="Installation">Installation</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="preparing-to-install.html" title="Förbered installationen">Föregående</a><a class="nextlinks-next" href="installing-upgrading.html" title="Uppgradera">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Installera från CD</h1></div>
<div class="region">
<div class="contents">
<p class="para">
	  The basic steps to install Ubuntu Server Edition from CD are the same  as those for installing any operating system from CD.  Unlike
	  the <span class="em emphasis">Desktop Edition</span>, the <span class="em emphasis">Server Edition</span> does not include a graphical 
	  installation program.  The Server Edition uses a console menu based process instead.
	  </p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
	      <p class="para">
	      Download and burn the appropriate ISO file from the <a href="http://www.ubuntu.com/download/server/download" class="ulink" title="http://www.ubuntu.com/download/server/download">
	      Ubuntu web site</a>.
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">Starta systemet från CDROM-enheten.</p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">
	      At the boot prompt you will be asked to select a language.
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">
	      From the main boot menu there are some additional options to install Ubuntu Server Edition.  You can install a
          basic Ubuntu Server, check the CD-ROM for defects, check the system's RAM, boot from first hard disk, or
          rescue a broken system. The rest of this section will cover the basic Ubuntu Server install.
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">
	      The installer asks which language it should use.
          Afterwards, you are asked to select your location.
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">
	      Next, the installation process begins by asking for your keyboard layout. You can ask the installer to
          attempt auto-detecting it, or you can select it manually from a list.
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">Installeraren undersöker därefter din maskinvarukonfiguration och konfigurerar nätverksinställningarna med hjälp av DHCP. Om du inte vill använda DHCP väljer du vid nästa fönster att "Gå tillbaka" och du får nu möjlighet att "Konfigurera nätverket manuellt".</p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">
	      Next, the installer asks for the system's hostname. 
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">
	      A new user is set up; this user will have <span class="em emphasis">root</span> access
	      through the <span class="app application">sudo</span> utility.
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">
          After the user settings have been completed, you will be asked if you want to encrypt your 
          <span class="file filename">home</span> directory. 
	      </p>
	    </li>
<li class="list itemizedlist">
              <p class="para">
              Next, the installer asks for the system's Time Zone.
              </p>
            </li>
<li class="list itemizedlist">
	      <p class="para">
	      You can then choose from several options to configure the hard drive layout. Afterwards you are asked 
          which disk to install to. You may get confirmation prompts before rewriting the partition table or setting up
          LVM depending on disk layout. If you choose LVM, you will be asked for the size of the root logical volume.
          For advanced disk options see <a class="xref" href="advanced-installation.html" title="Avancerad installation">Avancerad installation</a>.
	      </p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">Ubuntu:s grundsystem är nu installerat.</p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">Nästa steg i installationsprocessen är att bestämma hur du vill uppdatera systemet. Det finns tre alternativ</p>
                <div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
                    <p class="para"><span class="em emphasis">No automatic updates</span>: detta kräver att administratören loggar in på maskinen och installerar uppdateringar.</p>
                  </li>
<li class="list itemizedlist">
                    <p class="para">
                    <span class="em emphasis">Install security updates automatically</span>: this will install the 
                    <span class="app application">unattended-upgrades</span> package, which will install security updates without the intervention
                    of an administrator.  For more details see <a class="xref" href="automatic-updates.html" title="Automatiska uppdateringar">Automatiska uppdateringar</a>.
                    </p>
                  </li>
<li class="list itemizedlist">
                    <p class="para">
                    <span class="em emphasis">Manage the system with Landscape</span>: Landscape is a paid service provided
                    by Canonical to help manage your Ubuntu machines.  See the 
                    <a href="http://landscape.canonical.com/" class="ulink" title="http://landscape.canonical.com/">Landscape</a> site for details.
                    </p>
                  </li>
</ul></div>
	    </li>
<li class="list itemizedlist">
	      <p class="para">Du har nu valmöjligheten att installera eller inte installera ytterligare paketfunktioner. För detaljer se <a class="xref" href="installing-from-cd.html#install-tasks" title="Paketuppgifter">Paketuppgifter</a>. Dessutom finns det ett alternativ för att starta <span class="app application">aptitude</span> för att välja särskilda paket att installera. För mer information se <a class="xref" href="aptitude.html" title="Aptitude">Aptitude</a>.</p>
	    </li>
<li class="list itemizedlist">
	      <p class="para">Det sista steget innan omstart är att ställa in klockan till UTC.</p>
	    </li>
</ul></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
	    <p class="para">Om du vid något tillfälle under installationen inte är nöjd med standardinställningen, använd funktionen "Gå tillbaka" vid någon prompt för att komma till en detaljerad installationsmeny, som tillåter dig att modifiera inställningarna.</p>
	  </div></div></div></div>
<p class="para">Om du vid något tillfälle under installationen vill läsa hjälptexten som tillhandahålls av installtionssystemet. För att göra detta, tryck på F1.</p>
<p class="para">
	  Once again, for detailed instructions see the <a href="https://help.ubuntu.com/14.04/installation-guide/" class="ulink" title="https://help.ubuntu.com/14.04/installation-guide/">
	  Ubuntu Installation Guide</a>.
	  </p>
</div>
<div class="links sectionlinks" role="navigation"><ul><li class="links"><a class="xref" href="installing-from-cd.html#install-tasks" title="Paketuppgifter">Paketuppgifter</a></li></ul></div>
<div class="sect2 sect" id="install-tasks"><div class="inner">
<div class="hgroup"><h2 class="title">Paketuppgifter</h2></div>
<div class="region"><div class="contents">
<p class="para">Under installationen av Server Edition kan du välja att installera ytterligare paket från CDn. Paketen är grupperade efter tjänsten de tillhandahåller.</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
	        <p class="para">DNS-server: Väljer BIND DNS-server och dess dokumentation.</p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">LAMP-server: Välj en färdiggjord Linux/Apache/MySQL/PHP-server.</p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">
		Mail server: This task selects a variety of packages useful for a general purpose mail  server system.
	        </p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">OpenSSH-server: Väljer paket som är nödvändigt för en OpenSSH-server.</p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">Databasen PostgreSQL: Det här alternativet väljer klient och server-paket för databasen PostgreSQL.</p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">Skrivarserver: Det här alternativet sätter upp ditt system till en skrivarserver.</p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">Samba-filserver: Det här alternativet sätter upp ditt system till en Samba filserver, vilket är speciellt användbart i nätverk med både Windows- och Linux-system.</p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">
		Tomcat Java server: Installs Apache Tomcat and needed dependencies.
	        </p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">
		Virtual Machine host: Includes packages needed to run KVM virtual machines.
	        </p>
	      </li>
<li class="list itemizedlist">
	        <p class="para">
        Manually select packages: Executes <span class="app application">aptitude</span> allowing you to individually select packages.
	        </p>
	      </li>
</ul></div>
<p class="para">
	    Installing the package groups is accomplished using the <span class="app application">tasksel</span> utility.  
	    One of the important differences between Ubuntu (or Debian) and other GNU/Linux distribution is that, when 
            installed, a package is also configured to reasonable defaults, eventually prompting you for additional required 
            information. Likewise, when installing a task, the packages are not only installed, but also configured to provided
            a fully integrated service.
	    </p>
<p class="para">När installationsprocessen är klar kan du se en lista på tillgängliga tjänster genom att ange följande från en terminalprompt:</p>
<div class="screen"><pre class="contents "><span class="cmd command">tasksel --list-tasks</span>
</pre></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
	      <p class="para">Resultatet kommer lista paketfunktioner från andra Ubuntu-baserade distributioner såsom Kubuntu och Xubuntu. Notera också att du själv kan anropa kommandot <span class="cmd command">tasksel</span>, vilket kommer visa en meny med de olika tjänster som är tillgängliga.</p>
	    </div></div></div></div>
<p class="para">Du kan visa en lista med vilka paket som installeras med varje tjänst genom att använda alternativet <span class="em emphasis">--task-packages</span>. Till exempel, för att lista vilka paket som installerats med tjänsten <span class="em emphasis">DNS Server</span> skriv följande:</p>
<div class="screen"><pre class="contents "><span class="cmd command">tasksel --task-packages dns-server</span>
</pre></div>
<p class="para">Utdatan från kommandot borde lista:</p>
<div class="code"><pre class="contents ">bind9-doc 
bind9utils 
bind9
</pre></div>
<p class="para">
	    If you did not install one of the tasks during the installation process, but for example you decide to make your new LAMP server 
	    a DNS server as well, simply insert the installation CD and from a terminal:
	    </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo tasksel install dns-server</span>
</pre></div>
</div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="preparing-to-install.html" title="Förbered installationen">Föregående</a><a class="nextlinks-next" href="installing-upgrading.html" title="Uppgradera">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
