<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Wireless network troubleshooter</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a> » <a class="trail" href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks"><a class="nextlinks-prev" href="net-wireless-troubleshooting-hardware-check.html" title="Wireless connection troubleshooter">Föregående</a></div>
<div class="hgroup">
<h1 class="title"><span class="title">Wireless network troubleshooter</span></h1>
<h2 class="subtitle"><span class="subtitle">Make sure that working device drivers are installed</span></h2>
</div>
<div class="region">
<div class="contents">
<p class="p">In this step you can check to see if you can get working device drivers for your wireless adapter. A <span class="em">device driver</span> is a piece of software which tells the computer how to make a hardware device work properly. Even though the wireless adapter has been recognized by the computer, it may not have drivers which work very well. You may be able to find different drivers for the wireless adapter which do work. Try some of the options below:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list">
<p class="p">Check to see if your wireless adapter is on a list of supported devices</p>
<p class="p">Most Linux distributions keep a list of wireless devices that they have support for. Sometimes, these lists provide extra information on how to get the drivers for certain adapters working properly. Go to the list for your distribution (for example, <span class="link"><a href="https://help.ubuntu.com/community/WifiDocs/WirelessCardsSupported" title="https://help.ubuntu.com/community/WifiDocs/WirelessCardsSupported">Ubuntu</a></span>, <span class="link"><a href="http://linuxwireless.org/en/users/Drivers" title="http://linuxwireless.org/en/users/Drivers">Fedora</a></span> or <span class="link"><a href="http://en.opensuse.org/HCL:Network_(Wireless)" title="http://en.opensuse.org/HCL:Network_(Wireless)">openSuSE</a></span>) and see if your make and model of wireless adapter is listed. You may be able to use some of the information there to get your wireless drivers working.</p>
</li>
<li class="list">
<p class="p">Look for additional open or proprietary drivers</p>
<p class="p">Although Ubuntu includes support for a large amount of devices, some drivers need to be installed separately.
  Use the <span class="gui">Additional Drivers</span> tool to check for these extra open or <span class="link"><a href="hardware-driver-proprietary.html" title="Vad är slutna drivrutiner?">proprietary</a></span> drivers.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">
        Click the button at the far right side of the menu bar and select <span class="gui">System Settings</span>.
    </p></li>
<li class="steps"><p class="p">
        In the System section, click <span class="gui">Software Sources</span>.
    </p></li>
<li class="steps"><p class="p">
        Switch to the <span class="gui">Additional Drivers</span> tab.
    </p></li>
</ol></div></div></div>
</li>
<li class="list">
<p class="p">Use the Windows drivers for your adapter</p>
<p class="p">In general, you cannot use a device driver designed for one operating system (like Windows) on another operating system (like Linux). This is because they have different ways of handling devices. For wireless adapters, however, you can install a compatibility layer called <span class="em">NDISwrapper</span> which lets you use some Windows wireless drivers on Linux. This is useful because wireless adapters almost always have Windows drivers available for them, whereas Linux drivers are sometimes not available. You can learn more about how to use NDISwrapper <span class="link"><a href="http://sourceforge.net/apps/mediawiki/ndiswrapper/index.php?title=Main_Page" title="http://sourceforge.net/apps/mediawiki/ndiswrapper/index.php?title=Main_Page">here</a></span>. Note that not all wireless drivers can be used through NDISwrapper.</p>
<p class="p">Full information on ndiswrapper kept on
        <span class="link"><a href="https://help.ubuntu.com/community/WifiDocs/Driver/Ndiswrapper" title="https://help.ubuntu.com/community/WifiDocs/Driver/Ndiswrapper">this page</a></span>
        including troubleshooting help specific to ndiswrapper.</p>
</li>
</ul></div></div></div>
<div class="links serieslinks"><div class="inner"><div class="region"><ul>
<li class="links"><a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a></li>
<li class="links"><a href="net-wireless-troubleshooting-initial-check.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a></li>
<li class="links"><a href="net-wireless-troubleshooting-hardware-info.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a></li>
<li class="links"><a href="net-wireless-troubleshooting-hardware-check.html" title="Wireless connection troubleshooter">Wireless connection troubleshooter</a></li>
<li class="links">Wireless network troubleshooter</li>
</ul></div></div></div>
</div>
<div class="links nextlinks"><a class="nextlinks-prev" href="net-wireless-troubleshooting-hardware-check.html" title="Wireless connection troubleshooter">Föregående</a></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Wireless network troubleshooter</a><span class="desc"> — Identify and fix problems with wireless connections</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
