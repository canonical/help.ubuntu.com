<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vad betyder de olika formerna och färgerna på Startarens ikoner?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="unity-launcher-intro.html" title="Använda programstartaren">Använda programstartaren</a> › <a class="trail" href="unity-launcher-intro.html#launcher-using" title="Använda Startaren">Använda Startaren</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Vad betyder de olika formerna och färgerna på Startarens ikoner?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">När du startar ett program kommer ikonen på Programstartaren pulsera för att upplysa dig om att Ubuntu startar ditt program. Detta är bra eftersom vissa program startar omedelbart medan andra kan ta någon minut att ladda.</p>
<p class="p">När programmet har startats kommer små <span class="em">vita trianglar</span> att visas till vänster och höger om rutan på Programstartaren. Ytterligare trianglar visas till vänster om rutan när fler än ett fönster är öppna för samma program (dvs. två trianglar innebär att du har två fönster från samma program öppna). Om du har tre eller fler fönster från samma program kommer tre trianglar visas.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Program som inte används har genomskinliga ikonrutor på Programstartaren. När ett program kör fylls ikonrutan med färg.</p></div></div></div></div>
</div>
<div id="launcher-notifications" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Aviseringar</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Om ett program vill ha din uppmärksamhet (som vid en avslutad nedladdning) kommer ikonen på Startaren hoppa och skimra, och den vita triangeln blir <span class="em">blå</span>. Klicka på Startarikonen för att bekräfta aviseringen.</p>
<p class="p">Program kan också visa en <span class="em">siffra</span> i Programstartarikonen. Meddelandeprogram använder siffran för att visa dig hur många olästa meddelanden du har. <span class="gui">Uppdateraren</span> använder siffran för att visa dig hur många uppdateringar som finns att hämta.</p>
<p class="p">Slutligen, program kan också använda ett <span class="em">förloppsfält</span> för att visa dig hur lång tid en process tar utan att du behöver se programmets fönster.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="unity-launcher-intro.html#launcher-using" title="Använda Startaren">Använda Startaren</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
