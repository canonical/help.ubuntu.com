<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Mus &amp; styrplatta</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 18.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 18.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Mus &amp; styrplatta</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="mouse-sensitivity.html.sv" title="Justera hastigheten för musen och styrplattan"><span class="title">Justera hastigheten för musen och styrplattan</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra hur snabbt markören flyttar sig när du använder din mus eller styrplatta.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="mouse-lefthanded.html.sv" title="Använd din mus med vänster hand"><span class="title">Använd din mus med vänster hand</span><span class="linkdiv-dash"> — </span><span class="desc">Kasta om vänster och höger musknappar i musinställningarna.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="mouse-doubleclick.html.sv" title="Justera hastigheten för dubbelklick"><span class="title">Justera hastigheten för dubbelklick</span><span class="linkdiv-dash"> — </span><span class="desc">Styr hur snabbt du behöver trycka på musknappen en andra gång för att dubbelklicka.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="mouse-mousekeys.html.sv" title="Klicka och flytta muspekaren med det numeriska tangentbordet"><span class="title">Klicka och flytta muspekaren med det numeriska tangentbordet</span><span class="linkdiv-dash"> — </span><span class="desc">Aktivera mustangenter för att styra musen med det numeriska tangentbordet.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="mouse-touchpad-click.html.sv" title="Klicka, dra eller rulla med styrplattan"><span class="title">Klicka, dra eller rulla med styrplattan</span><span class="linkdiv-dash"> — </span><span class="desc">Klicka, dra eller rulla via tryckningar och gester på din styrplatta.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="a11y-right-click.html.sv" title="Simulera ett högerklick"><span class="title">Simulera ett högerklick</span><span class="linkdiv-dash"> — </span><span class="desc">Tryck och håll kvar vänstra musknappen för att högerklicka.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="a11y-dwellclick.html.sv" title="Simulera klick genom att sväva ovanför"><span class="title">Simulera klick genom att sväva ovanför</span><span class="linkdiv-dash"> — </span><span class="desc">Funktionen <span class="gui">Uppehållsklick</span> (svävningsklick) låter dig klicka genom att hålla muspekaren stilla.</span></a></div>
</div>
</div></div></div></div>
<div id="problems" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Vanliga problem</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="mouse-wakeup.html.sv" title="Musen reagerar med fördröjning innan den börjar fungera"><span class="title">Musen reagerar med fördröjning innan den börjar fungera</span><span class="linkdiv-dash"> — </span><span class="desc">Om du måste skaka eller klicka med musen innan den svarar.</span></a></div></div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="mouse-problem-notmoving.html.sv" title="Muspekaren rör sig inte"><span class="title">Muspekaren rör sig inte</span><span class="linkdiv-dash"> — </span><span class="desc">Hur du kontrollerar varför din mus inte fungerar.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="tips" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Tips</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="mouse-middleclick.html.sv" title="Mittenklick"><span class="title">Mittenklick</span><span class="linkdiv-dash"> — </span><span class="desc">Använd mittenknappen för att öppna program, öppna flikar med mera.</span></a></div></div>
<div class="links-twocolumn"></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html.sv" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html.sv" title="Mus &amp; styrplatta">mus &amp; styrplatta</a></span>, <span class="link"><a href="prefs-display.html.sv" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html.sv" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html.sv" title="Användarkonton">användarkonton</a></span>…</span>
</li>
<li class="links ">
<a href="hardware.html.sv" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a><span class="desc"> — <span class="link"><a href="hardware.html.sv#problems" title="Vanliga problem">Hårdvaruproblem</a></span>, <span class="link"><a href="printing.html.sv" title="Utskrifter">skrivare</a></span>, <span class="link"><a href="power.html.sv" title="Ström och batteri">ströminställningar</a></span>, <span class="link"><a href="color.html.sv" title="Färghantering">färghantering</a></span>, <span class="link"><a href="bluetooth.html.sv" title="Bluetooth">Bluetooth</a></span>, <span class="link"><a href="disk.html.sv" title="Diskar och lagring">diskar</a></span>…</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
