<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Install the Flash plug-in</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-browser.html" title="Webbläsare">Webbläsare</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Install the Flash plug-in</span></h1></div>
<div class="region">
<div class="contents">
<p class="p"><span class="app">Flash</span> is a <span class="em">plug-in</span> for your web browser that allows you to watch videos and use interactive web pages on some websites. Some websites won't work without Flash.</p>
<p class="p">If you do not have Flash installed, you will probably see a message telling you so when you visit a website that needs it. Flash is available as a free (but not open-source) download for most web browsers.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">How to install Flash</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Click <span class="link"><a href="https://apps.ubuntu.com/cat/applications/flashplugin-installer" title="https://apps.ubuntu.com/cat/applications/flashplugin-installer">this link</a></span> to launch the <span class="app">Software Center</span>.</p></li>
<li class="steps"><p class="p">Read the information and reviews to make sure you want to install Flash.</p></li>
<li class="steps"><p class="p">If you choose to install Flash, click <span class="gui">Install</span> from the Software Center window.</p></li>
<li class="steps"><p class="p">If you have any web browser windows open, close them and then re-open them. The web browser should detect that Flash is installed when you open it again, and you should now be able to view websites using Flash.</p></li>
</ol></div>
</div></div>
</div>
<div id="alternatives" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Open-source alternatives to Flash</span></h2></div>
<div class="region"><div class="contents">
<p class="p">A handful of free, open-source alternatives to Flash are available. These tend to work better than the Flash plug-in in some ways (for example, by handling sound playback better), but worse in others (for example, by not being able to display some of the more complicated Flash pages on the web).</p>
<p class="p">You might like to try one of these if you are dissatisfied with the Flash player, or if you would like to use as much open-source software as possible on your computer. Here are a few of the options:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p"><span class="link"><a href="https://apps.ubuntu.com/cat/applications/browser-plugin-gnash" title="https://apps.ubuntu.com/cat/applications/browser-plugin-gnash">Gnash</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="https://apps.ubuntu.com/cat/applications/browser-plugin-lightspark" title="https://apps.ubuntu.com/cat/applications/browser-plugin-lightspark">LightSpark</a></span></p></li>
</ul></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-browser.html" title="Webbläsare">Webbläsare</a><span class="desc"> — <span class="link"><a href="net-default-browser.html" title="Change which web browser websites are opened in">Ändra förvald webbläsare</a></span>, <span class="link"><a href="net-install-flash.html" title="Install the Flash plug-in">installera Flash</a></span>, <span class="link"><a href="net-install-java-plugin.html" title="Install the Java browser plug-in">installera java-insticksprogrammet</a></span>, <span class="link"><a href="net-install-moonlight.html" title="Install the Silverlight plug-in">stöd för Silverlight</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
