<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Flytta ett fönster till en annan arbetsyta</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord</a> › <a class="trail" href="shell-overview.html#apps" title="Program och fönster">Program och fönster</a> » <a class="trail" href="shell-windows.html" title="Fönster och arbetsytor">Fönster och arbetsytor</a> › <a class="trail" href="shell-windows.html#working-with-workspaces" title="Arbeta med arbetsytor">Arbetsytor</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Flytta ett fönster till en annan arbetsyta</span></h1></div>
<div class="region">
<div class="contents">
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Se <span class="link"><a href="shell-workspaces.html" title="Vad är en arbetsyta, och vad har jag för nytta av den?">Vad är en arbetsyta, och vad har jag för nytta av den?</a></span> för information om hur du aktiverar arbetsytor.</p></div></div></div></div>
<p class="p">Använda musen:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna <span class="link"><a href="unity-launcher-intro.html" title="Använda programstartaren">Programstartaren</a></span> och klicka på <span class="gui">arbetsyteväxlarknappen</span> nära botten.</p></li>
<li class="steps"><p class="p">Dra fönstret till den arbetsyta där du vill ha det.</p></li>
</ol></div></div></div>
<p class="p">Använda tangentbordet:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Välj fönstret du vill flytta.</p></li>
<li class="steps"><p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>→</kbd></span></span> för att flytta fönstret till en arbetsyta som ligger till höger om den aktuella arbetsytan på <span class="gui">arbetsyteväxlaren</span>.</p></li>
<li class="steps"><p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>←</kbd></span></span> för att flytta fönstret till en arbetsyta som ligger till vänster om den aktuella arbetsytan på <span class="gui">arbetsyteväxlaren</span>.</p></li>
<li class="steps"><p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>↓</kbd></span></span> för att flytta fönstret till en arbetsyta som ligger nedanför den aktuella arbetsytan på <span class="gui">arbetsyteväxlaren</span>.</p></li>
<li class="steps"><p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>↑</kbd></span></span> för att flytta fönstret till en arbetsyta som ligger ovanför den aktuella arbetsytan på <span class="gui">arbetsyteväxlaren</span>.</p></li>
</ol></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-windows.html#working-with-workspaces" title="Arbeta med arbetsytor">Arbeta med arbetsytor</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-workspaces.html" title="Vad är en arbetsyta, och vad har jag för nytta av den?">Vad är en arbetsyta, och vad har jag för nytta av den?</a><span class="desc"> — Arbetsytor är ett sätt att gruppera fönster på ditt skrivbord.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
