<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Användarkonton</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Användarkonton</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Each person that uses the computer should have a different user account.
 This allows them to keep their files separate from yours and to choose their
 own settings. It's also more secure. You can only access a different user
 account if you know the password.</p></div>
<div id="manage" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Hantera användarkonton</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-add.html" title="Add a new user account"><span class="title">Add a new user account</span><span class="linkdiv-dash"> — </span><span class="desc">Add new users so that other people can log in to the computer.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-changepicture.html" title="Change your login screen photo"><span class="title">Change your login screen photo</span><span class="linkdiv-dash"> — </span><span class="desc">Add your photo to the login and user screens.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-delete.html" title="Delete a user account"><span class="title">Delete a user account</span><span class="linkdiv-dash"> — </span><span class="desc">Remove users that no longer use your computer.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-guest-session.html" title="Launch a restricted guest session"><span class="title">Launch a restricted guest session</span><span class="linkdiv-dash"> — </span><span class="desc">Let a friend or colleague borrow your computer in a secure manner.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="passwords" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Lösenord</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-forgottenpassword.html" title="I forgot my password!"><span class="title">I forgot my password!</span><span class="linkdiv-dash"> — </span><span class="desc">Advanced techniques for resetting your password</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-changepassword.html" title="Välj ditt lösenord"><span class="title">Välj ditt lösenord</span><span class="linkdiv-dash"> — </span><span class="desc">Keep your account secure by changing your password often
    in your account settings.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="user-goodpassword.html" title="Välj ett säkert lösenord"><span class="title">Välj ett säkert lösenord</span><span class="linkdiv-dash"> — </span><span class="desc">
      Use longer, more complicated passwords.
    </span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="privileges" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">User privileges</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-admin-change.html" title="Change who has administrative privileges"><span class="title">Change who has administrative privileges</span><span class="linkdiv-dash"> — </span><span class="desc">You can change which users are allowed to make changes to the system
 by giving them administrative privileges.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-admin-explain.html" title="How do administrative privileges work?"><span class="title">How do administrative privileges work?</span><span class="linkdiv-dash"> — </span><span class="desc">You need admin privileges to change important parts of your system.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="user-admin-problems.html" title="Problems caused by administrative restrictions"><span class="title">Problems caused by administrative restrictions</span><span class="linkdiv-dash"> — </span><span class="desc">You can only do some things, like installing applications, if you have admin privileges.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html" title="Användarkonton">användarkonton</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
