�PNG

   IHDR  �  L   
U��  zTXtRaw profile type exif  xڭ�Yv��D�1��f8hת��kHQ�e[��'�"�D"��ĉ  ������r���T*o��+��|�M���q:������ϫ���8m��<����m����:�����|�{k�����y��?��y}|�>�������{<ٮ�ώ��(>~���V˧���|r|^���c(>��J�g����x_��{.�L�nG�a�ׅ��ߚz��wp��3�e�:���.D��.��χ�-�d��=������6�6���O�ey��j��k�ׯq�_W?]�{���k5??��j�����.�u��Ax=�|r��'������l����zE�[��ަr��nȊ���w����7�n|W��$���d��}s��r����t�!F�}���i|�+Nj~Ą���Y���P�5w��㦫v�M��3w#�_~��6<G�䜭;��+8�u�_/4�#�<����߾�~ɯ�k������H�=��ut�a������g��G'��م�2#*��0d�A�����.%���!d�Cv�l�)�6��?.��$mH!��o�b�c"~J��PO!ŔRN%��R�!+�r.Y��K(���K)ՔVz5�Ts-��V{�- ߩ�����z硝�;ww�>�#�4�(��fF��ό3�<ˬ�;�
�_y�UW[}�M(��λ���P;�ēN>Ŝz��/��g�~��^sO���)5,/�q���.��$�gx�G��^�c�|f����s����H�A&9g9y��|:�廧�V���͔z���S����o�ym�J��Gʨ6�}��ub�Q�d�ؠS�i�����y�d �j���yrs#Oyʃm�����Xu��
7`���ڻ�=f-����lq%�0ڊ��P.�Ƕv�L�Z�W�����>��5���1�d�@ڥ��Ƀ6������&y�L۽
ͪM��n#)�z���� ��exϦwZU��5B�oߏ��*Ԫ���-�2����;�X�~l�X�[�܇�u����iK
c�u�������~'v�#��&�3��ѳ�j���yX�OV�ń�����_|����aC��g�_��w����b���/�ڀ��לu�]��L��X~��<�ԁ��II�ˮԆ�M ���}G�B[9ө�i��}��μ��5�c�\%m��,�]P@!��R_a��f.��U��`6��2��`��|(b����$M�Їs�'���k��_��̷�k�Us��b<�y`�JQ���5=��
�֯�\��ZegPq`��v�Ӧ�������r�<�5�3h �P�<p���ka������u0�s�V�0�И�vg�����:b�r8#�J�Gv'a�<\��P� W:�f�ɹ&q,���H���)�=T��<6o*E��,��1'��!V��AΰW��?G���U�Go��FH�S~����:�j_���da=q@��Z�2��v���:\9�����t�XFjY��F1T��3�6C-ͧ�>3���k�z����{�CJz
ⴌ���+�`�� ���U�G�B�g\��tg]f"��,$۫Y|� ؃P�9�]29I�-�BT��J#R|��(]e�RL,b�����r�d;��#O2��[�
�5�ڎ�&_Pw�E~��B�;��R��lY;�~'̐8!e�Y�|��,��U|a��7v�J��~����X0�
�ިC=m,1"2��k���}'��+^f[�bs�_ۘ/�v ;]�#�G��Z�a���|��11�N�xQ��U���d��dRh��w:�8� %��Ŭ�&"������Ö����s��c$����f��d��R��q�(�.a�0�@���J�] ��K�0�u@�5-�I�����s`��yH�f�eV�!�#y�0~���ݞ���H��5oO��jNq;ֺ�P�.X�n���`�}�(BNQT ��Z���A�.�z0��k���ԏ��=��e��_b���b�
�(g��ש��	bkD ��!��1�IQW'uj����gv��^M�)� Ɉ�^�� �͡'���F�R�|MЅ�&����g'�PHHi��ܕ���AP�S�*	��j:"g	�Iwбs9TÉ)Nܙ���@� ����,�ZO�V�j2e�w)� G4a�0W�u�Ax_[�ӧ��K��	�R����<�LG��,V�Y�����s�����!`[΢���S?�	Q#��A�p���# r{k��6u�2s�zs���\HZk��+cc���^qD�B!��!�X�%��<^/CN�_��.*!4���i�ꌪ.1H�Y9�مꚔ��E�kH�����Er����$�$���y	*���vwR�nG!i�"���=�"�d_����ug�A�� 6S�wC�ݲZ��	�EH* &&,Ш�Q�>C�S�#-�)+�Z��v-y4Ȉ���
��X�AJy��_��e�s�^zD��e ��Ix�y(<��P�{��ɕN��omfI�z�W��B$��	�?z}�	C������JT��&M���n��bT�LZu�
�y�Ax�Q΄=MԼ��;r��P	/�P���I9�d �e�UB����&� c��"s�}G���T���+�����LF��J��D� �.�S��G��5��T
�������"<�R@ʬ2%M'XGJ=Ȗi0
w"9`Z��+S9$H�K-����@@����+Q�5�@;)َ|m���=�*���}��"�5^�:�<T ۈ�T&`��MԒ����0�Vʸ�U�w��1Cn[[z���z��Ыs�;ʦ���F��hZ�(����H�Fܩ3�1���3��G8�܂�Ub���~4�];��ƴ�/��i�!�C�O!�m�W����v��;Bʠ�� �����\���@�9���f*R�G�n��0S�M�ͷ��=��$�\H�5U"�?$0P���b��޵F$lÅ�N��RNy��$�!�B�7���Y�E�5H����1[҃Ȉ}��{JZQ�JZ����)��д�ג`MG)p����X	V����ikI2RkV�;�ӌ�ϸ0�Ɵ@n�9\&̶ӜIIۆG��t_�����{��F����3펽ɀ���5�6w��E�����r�:�����F�i�*�P}�-�'��eN?��r��M1v"���T�J6��1}���gY1�;]팛`Ha��O(���O��-�x�y<3���H@(ѳ&Pɣ�ݟ�z1AE���xe3s����>�m�|�?�OiQ�n���2��J�%��uO��Zq�"<R��@]�gx㴇���J�~[�nҿ���d�8P9E�����2Г�$1�Ev�D�-�EV����S���� ��Z�n�mW��G�2�	i�n9�@it=��&����`D����A����D7A��ɍ6���4�O�����t��z��z"�ߦX�c4յ���w�Z�>z�b��.��5���kQkOT�5�M[����k`8�2�VB0��XJ�B�B��̽����~-��*IL�7�t�Zu�ΩN^l�AUf����7���=�,�O���3Uj�T��Z�&��3�E�\#3���:[��3�w��M͋��N��.l�^�7����� ���i]����.?U���Lݰ�W7��&���HI8������V����Gk�i�=D�*�D����-a����C�"��]GP(iq_���@��/k��T�1ĕ������f�g�Zf�Q�r~7� �W�����;�L
Y?�[ $�;��)E+���Q	y�\hsD'j0Č�$ݎw�!�����K��l�RU�|�j@|V�t���:l��)ԅ>A�i_ig[���&�r�L��z�o�',?�+���g|���ܜv���$8�\BՓ�Z��.0�[H)��J#c��&�Z'�6r4"�@lP�H�L��;�k�B.F�IqХy�	̓,������� ->��Q9��(I 7��d�)nڪ��Q�&<�</�؇����l��T��^�R4@ygkA	�l0���B�z�j�p����U<Ҍ�8�j.vH�'����
7��?U���ޓ�����7!SUw�I�q9����][d`&h�Y��AT��W-�Q�:�����En��'w�W$��=B5~Ϩ���t��ά�O2'��!��dL�ؙZ�ָH�e�<�V�l�{㮕�!�^���=����m//r���t�
5�s�w�J��#�vR4P�ݳ�G
7��`�
��!e�=���� ��`��<u�AЇO���]rG���O��!���l���1�_�L�1Y�J?��F9mh1��`@x�(��/��j!a)�S���(�Ɉcb:Y无u:trwՠ�GO ;�y?8W��֙����Zg��b�o
��D6�+�� �z�h������z/iy8�H�3��!���&�
��L~9�P���W WZ����R������I���u�h�����_lظ����h�z7~����_���A(���٠�8P��Ϡ�!��a���Y�E����6�u�S�T%=\��r��l@�K������o��¢dڶ�!�=S�h[ �&yu@u����`�q�|B<1S�vA��V�_��Xh�9��'h?A]-͐�=]RJ�G�[P�BPS0EV�F{S7YJ�w�.K��!����x����v��1I���NŲ ��ͭ1���9)l����]Jk���T[��d#���bl�(K7�5��eԢ�5��[�ϩP?��J��ynB�Jl<�
��d-6��-����mp�i��X�9d�h8
B�O�
mQ�Rr��*��1��I\}�$�|TQ`v�ck�W[��s���7��%Ή1l\uhp.3+a�$��h�t g�*L�����e����q� :��\�qC+�t�%G��gI�,��?]Y��T�u�&%�(|ELt$�V�\��G���q� �U��:��,~毫Vo���A	s�'�>2uʡ]�M�W��C
(-��¾"��m� �H�ں.�U�~ }���(S5+;
�rgb����Q�=K�;�Q=����Fw+�c����3~�.h=���^M;_*Oڐ�j߹Q��q� ����Z[�"��!%�Jq!Vf��A�,󘒚0J�h���;q�U�o%k���<CR��R=h�FM�������?����6;n��,�cj�A��	P8���%�1 �.�;�uvJ�>"���c�%;wE�F�E��dD�����cu�$��:2�����p������Q���{S���"&���3��h1�ƤH\N���������y�G�i�X�跊 �!��Ȃ:H ���ǧ�>Sg�J�"���FAJ��r��m����87�vI�4r�Vg>)�𑐑P��XI���H����)
 �c=�;/�j�;@$ZMM���(�y� 	]��<@_�3xQd���\�!�q��n�Y	Q��$����#�B�m����Ø}���,�OB�R@���%Ġ��ٔޚ�Hb 8���[�@/`�K�TX1Ӿ�.��Ukh�qM�2G�c�yY����]��VD�t�y������U� 
�"�2���]&6#��(��1
�^�� ���,n���Y�ŉ?bS�
(<!�`;ь�r����dPgia+���Ic���@t��:/��^���FthRZ��hy�I�V��2��v�:�g�(��o]&3mj�L�o�&I	��Нs�]��24� %�Vq�Ա�V��X� ��d�j�����֑��� ���a�M܃,o*Mn�Z��M�礿x����)��ܞMe�3>�m�����~|4�{��?9j�O\�c[����}�U'�>�i��dz^g!B���|5��O�b��s�����Y�$0Z3u�L'؂����g(���0��Q��L�[�yO�}A�m9�q���.��=1_��ᵧ!+`O�:� ^[m�1��ʳH,���j02<�����s�٠�8�_wP��jf��@���'��#�0�^ř�g���ɂ �h�VT��Z�����2��YkY+�	����"ڐ�^�vU�(��a� n?7.�`$a�]O�},�Y�%�Ѷ�縦U�5�\�c⁦l-Crw�"�@�-� �:6�A�J٣�ߠ���;�F��-�}5��m�ɴ�_C�~G�`wQ
>���Jǘ���[6��,
ӓ8���Fp1�ys��^Os�� ��z��\�>lhp2v�9*Fյv�� ;�*��<7�G1^��o���p��:b�C���Dv��(��s^�˷�}�9z�Zg�)ʡa2���
��
{7qt���i���ʍs�*��  �iCCPICC profile  x�}�=H�@�_[��f�P�,��8j�P!�
�:�\�M�G�����b���YWWA� qtrRt���Z�xp܏w�w�`��4�m�t�L�cb:�*v���0���,cN��_���.ʳ���9zԬŀ�H<��&� �޴���+�*�9�I$~�����A�)���<�@,�[XiaV05�)∪�L{�r�⬕*�qO��pV_Y�:�!ı�%H���"J��U'�B��c>�A�/�K!W�(C������w�Vnr�K
ǀ���:v�z�q���~���+��/׀�OҫM-r�m�MM�.w��'C6eW
��r��}S��׼��8} R�U�88F��������=���FUr�iV�  xiTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:61894402-3936-457e-83ae-3e0a4ae8daac"
   xmpMM:InstanceID="xmp.iid:29153034-9df1-4d4e-9916-74c6160dfa65"
   xmpMM:OriginalDocumentID="xmp.did:174b53ee-173d-4965-a4e7-2b3292ca8336"
   dc:Format="image/png"
   GIMP:API="2.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1663187550517887"
   GIMP:Version="2.10.32"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP 2.10"
   xmp:MetadataDate="2022:09:14T22:32:30+02:00"
   xmp:ModifyDate="2022:09:14T22:32:30+02:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:58f17fcc-49cc-49a8-9707-3f47b8e2a84a"
      stEvt:softwareAgent="Gimp 2.10 (Linux)"
      stEvt:when="2022-09-14T22:32:30+02:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>n8�   bKGD � � �����   	pHYs  .#  .#x�?v   tIME�	:��   tEXtComment Created with GIMPW�    IDATx���w���������~����ы�tD�*�Q<I,�&�$��@�X���؂5�XPc	#$�� +�J�*�
������ػ��z�E^��c�;�3�������}�;FiI�-  p\��X>�����4Bp�&�  ��apu>   ��t� (�4   |�   ����|   ���4ApuΘ   ���ɇ��1�   @r��q   5�W>��W����^:l����?���_�Z�a��q9��   ����E�.I�o�A�%%%�q�<���';��
e�����������(66���`�   �y.�K��v�6m�\��e|�3Ϛ�O>����Z�b�.��u�������_�R���Z��mޏ��b  �N�����A]C�-Ρ��-��o�7�������]dҸ�����C"�?%D�!��v�կJ���R��&�׵�cԫ�S�%�^_W���j r]8&J7N�������Ů�Vo�-�+�������}�i�ڵn߶l����?�IcǞ����V�kŊ���?Ȳ,M<�4��сB�mk�С�|�]����ȶmM�2���E�:  h�!�����������u�#Mݛ���;ˏ��yR�6�Խo�k�����
�~v�f���;Yy��D��[�˟?�'�W�����U�b|�xE�����2K?]���ظ��E�FÆm�km��'����y�7s��k������OS��}����O>m]���Ç���˲,]~��u�-��Y��[n���3Y����V~~~����L�  ������jǎ�m[]���+.פ��λ��Ǟ�ҥ�)2"�����W�В������×�U���=�?=5���LC�{V��XW��J[���7��顺nj����0���n=�q�Vl)��a����(�Lr*���G[������қu�� I�*�h�	��0�fO��,PN����}%���ڽ����Oג�K$I����yn=�^�$i{�K�	���h��Y��]�b#LE�~��X��lW��n�v�W�l�/~B�4i�4I�G.o���r�~�Q��j����B�عK�������9��@O����裏4u���s�ҥ*)-��cF���~^�qx�_y�eڸq���z�^[�DW^qy��Ѵm�T�<x������<\.�n��v�x�`=��3z���t��W+*2Z�-M�4Y�ij��~��|�]�7N��q-�g ]1!Z!�O��׫hz��Dm�W�K��Տ���_V����s�(�fZ�^ZY�����]�=�a=Bu�9�~ۚ<0Bn[?|2[g?�%�%��Q��VK����ңuO��;��J�rg�"BJ����k�[V�Nl���9]��]��Ϻ��"��7g�����;��m8�]秗�T����d���Q�$I[�|۪}V��_t�E~�:TÇ�{�.�$}���>Fz� ���"�딱c�֭�$�kj���."<L�&MԻﾫ�=S�����/��R��s��������٣����5{luL���0S����|���_L��_Vꝍ�����2���J�*��o�>T���y�u�Y��[�7~���}´��x��5<R't�#���H�2�W��;�W��.1�z���[|�P;r]
s:kH��Ǘ9����Vo��{�'O�֌u�6��+��h���M�?j�I�v��)�Vj�TI����Zu����d���'����z�N�U��o߾V��:�� @`���k�Yg�[nш�#4|�0M?^}���3s����ou��������)..N��r�1s�I��=+Aw���CŞf��H��7חꉋ���J}��B�l����P���N�E����x�~v|���'8u��;�{{���!�ȣ#���vq�(��yb�~wV��~#_�T�)�~�]����}��B�a�~zj�~Q����(�0�u{���jt�����8�� ������t��.��/���_��A���/t���?�:TݺuS�;���/׻ﾧ3O?C��8f��>05D�Q��(��uӐ>�5M�}R�g>.��������_��>�:�w������(��+KdVM�1w��:�Cjs�u���ҳGEi�������ݟeK�K,%E�o0)�[`��IT�!�G�p7��m����#�0�����n{j�w�����)Ӧ�=oH��Z��ԔTe�d7Z��_}-I�ݧ�l[:x�$)1)�Uǘ����;�k���:9!��u���)I�ѣG�FM�i<x���#Џ�}{���|@_|�^��2Ðf�5]����l٬�v��Κކ�u�u{+��gru�G�(�eK�>��W]��`��q�U%���^���7�ʾ#n�[�4 ��w�N�X�or�b�M��s7��<-Z�O�ռW�����X���S����e�۪�E�^���g4~3���Ct�Ē�c7{������^����7����4Z��/�"I:�3$���kop|�	������$I�/nr�E�IR�{Zw�&�y������>��٫g�]�M�lҡ�<m۶]k׮S��}�֛~�t������נշO����aNCSC405Da!��"��T]�XZikG���W��#ץ#%V�����uSb4�{��c�5D�{�iG�7\{,陏��12J�L�Q���Ltj��p�u��P���;ωW�.NI�]����,�������ߞ�+O�՟�*���k�.GG���D����7=N�SBt��H]rj����љY��Ԟ�GOn����Fjx�P����Ύ��#��ʢm7�9����є����O�z�����V������c�h�B}����G?�w���H�8�D�:�ٖ�7�|K�����֪c<����ի��sϽ��z�.xN_~�����4;#��?�N��M  TXD�v�ޭ��_�����ј1ct��W����SSS4b���z�����
����Jr�+�}�{&:5eP�,�m74*��ջ�7��G�*(��jg������)�W+�ģ���%�D�mI������2�m}��\�r�o�tQt��/wW�̂f��̡�r���3����wĭ>�#Iڸ�R���a]3)F##�_j���z�Ɛ�������+ܶ�8-Z)1U�m��s���9��7��9�mߜ����ƍ뼶aÆ:�j�z-q�5W+��!}X5�z���^�)-[��v�ڥ�ݺj��_|B���x���>���K���F]|х8p�$i�֭Z��EZ�f�L��M���ظ�V�q$/�� �qf����1?0;AK����h�{׆��=S��Q��+�/k�z-�r�t�ͷh��u�nk������;~�N�0�M�����#�>���/�������ݨI'�i?Nq5)   jj�|��m�q�!N��p�ݚw���nkڔɚV}��6�kʤI>t��������ڻo�$)�G�ƍ;U�7K���mޏ��   ��܊�z�6l�X�5���FdT���׿tʠ���x]��鲟���ڰ6�pnY ���YOU�hлW��A�;�  ��aPu>   Ӄ0�s1)   ��:�0�4   |�6gL   ��|�Q   �    �øꪫ��  Ǚ5=�Р�{��!�DP   �C_    �:    �:   p�rv���  ��LA��   �����Ύ+���0�5D�Κ��N�n�RԣGWEEE�  �{���L{�TVV�>��K���r}��7�����ގ�3�u��~t��g���%˲�<ޥ��'	  ����^�02MS[��֝w<�%Kޓm۵��A�?����S/���ƌ9In��`  ��i�r8������k׾f��v�߿��6Z�_��b���t   p�s8�*(,���ъ�j�t�#��H�2e���\ ɢ   ��MS���3�����E�a�A��K�>=���EH   �a��j���}�56�nx�p��>���B:   � ��(.6JϿ��PcӚ�2��y���3�$Ƥ   M�x�:��:��3����Z9����C�fS�z�N�7   h�4�s�~�4���Wj�۪u��?z�Iп!   hn��,�[#G���Ֆ����Y��"�   -bY�Νuz��^A�ք	�|w ��&33�F �!<�G'�ipy�{ԻwOm�bU    HKKQCa��A�[��$u   �El�V��]\��)�u   ��Iݛ�;*�   hu   ��   ��   �   �   �:    �:   @P   @P   @P   �    څ�&   �d���$��v˶m z�   �:   ��`�  A�4M��)��[�,�,���p:e�d۲,K��I�-����b�L�ûnնly�c�ܞ�!����ٖU�P�:uI��۪�=[�m�d(���4  ��p8���0$��eH��!���>�� n��=����@�̒-�0dȨ7TK���ա�W�$C�m{�e{O5Ojo�>z� ���Q  ��8�m���U��)�4�˨�]�CmVlC~�Y�<�Z��5�׻��_k5k�^O���{<IF���� ����}�Ys(�ey�0�����m����wC�m�z��m���*�_஽O۲d���}�b�@�5�xS�@P �XO��,k|�����0}�]�裺��y�G��x��X�%9
� �  |o��7LS��6k�o�E��!_�w[_p��K���:�Tj<�j\��Z��v�Ps< �:  �XN��T�7H;�!U��j�e�(����R5Ӌl�0�Z���>MS������!˲�N �V�}��mƩ.  ��x�=������3z<~s6?����0�g��q{��Y=��:��셯ޖ���n�4MY��ޑ75�'�{�Q{{ Z�u  ��eY~s����_nۖ�.�Vhn^��x<R�0]�۲��Z�uu�Ws�H�P�    LӐ�pzy�<���_,�Eu  �S@���� A  tbPo�ԏ ��Ť    A    A    �   h/\L
  ЁӔ���=����+�:  �L�3L��!��N��	v�C���s����
/!!���<��n�hw�iz�nkT�.��ki۲,��v7����>��;ֶvm���  �5f��ޚ�_;���f������t2MSOݓH�0�p:��a�4꾯��kK�����W � aK�e˶Z(�-_Kۖ]ߍ�����^�;m4�]m�����`F�:  A��͂ӔC-��m�7L�;��o�d�{����.�Q5��{�e[��_ϸ��m��v�j�BuO���s\�Ô�8���v��=�-��v�Ѻ��ےeydU�A�tT�\wYc̪6n�X;�m�����S��\�<u�Ű,���:��Y�FI���M�F����-k��Z�>�:  ��i�0�A��x�]+�Uo�!��-����*����0��Pg�G�0e������:�._�!�4\�ظh�t�>�����ڶ)�m��Mڶ��`�W5{�-���n��)��6��;f~��� �����o��զ����FȲ��x��xd����k�3۲|��>*k��s���uPs؂e��A���|��۽.�u�#��)��T{Y��4�>��?����u��Q�,����5֓�X�����z� 8�9�_ �x���}�A���W��������m�>:����P�:�Ͳ��w8��^��=l˒-�0���I��e۾aI��������Q}���c��v;ْ��>3�8����j��������}u  �.�������	"5�8��vȖ��U��	�5zEӐ�i��0�P�f��Z��?N��g��'�_�]k����%=��>�v;���nԾF���thOuk���u� @ݠ��r�续,�������2�	L��7�{K��6��]����{��ڵ��u�uOjZy:�䱪���C]��;����o4�����k���  ���)g#�W� �97>�m[n��7�0�ބ�fX�{�e5:F���T+�מݣ%1�]��O��c�c0��𪪓
���j���N6��kn����>�:  8�TϚ��5f�1T�A���%�n��Lb��x�Q�0k�p�� ڥ����c�1�f�1�������%�o����kO��kj��5�k���  �����d�	"��m�>z�g7F����/�4;T]�h���ҽe՜�&�)�����^�������"������G�f~퓆��#��_���}�W]����c𞘙uN���U��ڲ����{��mU}�kuۿ���#� ��7ì3�v�`W�-Y��Xm����u1]K{�n��O��-��_�ZyH۲��K^#`�=�-�^�a�fPo��:B}��c�ch��������ò�9CQk�@?��N'� �B�%�"kݙԮ���s��w��껙�M��Z�G�m4�n��a�l��N�QWG�ޔ������ԉ����ެ��wSA �����	��l�j�[m�z��������ls*mi]��`ۖ�.��p�P��km�ީ.����_G~m��ڲ���3�qgR   ��   ��   ��  :]{�����Q   �    �    A    A    �    �   u    u    u   ��   ��   �   �   �:    �:    �:   @P   @P   �    �    A    A    A    �    �   u    u   ��   ��   ��   � @{{��h���7ܨ�g�Я}=��Ξ�y�:  h�����/��h���4���~�UVV� �#�.x��u  ������i�;˲��x�۰��r� ���֯_��^~E�v�TiY�b���޳�~8{�ƍ;շ��￯7�xS����c�w�^��gk�ԩ�un��Fm��0@g�q��,]���<�LO׵�^�aÆ��k�ӎ�;}�9��Y������;��}��5g�\m޲E���g�/����#3z�~{�o����z�u��a4Hs��Q�n����>�H���?����Wgk�{֬s��_�t��A��/Q�~}���Ղ�We�K�\s5A  �[���D�����W�O����]yyyڲe��o���O?�����k��aC��0M�[�N<���֏~�C��n߱C���2d�*�˵c�N�v����gԧO�(//O�t A2Cݻwoվ��۫?�X�*/��'�~����j��=���Pii�֬Y�GyT?<��{z�JII�eY~u�������v��Ï<���$EGE�߯�^~Y��2��  ������WH�n��f���G�TQQ���"IRNN��,]*I�����g?��_�~��u�~���p�m?�أJKKӾ}��_^���J-~�U�t��`�sZ�x�$���+44���*++�zPÆ�o~3G[�m���{t�5����3��?�ײ>І�UYY��W�{yx������k��n��yх�����J͝��}�ٲ,K�eփ4�� B�aa4B�=�+55U��ٺ��k���=5l�0͞}�$i˷���˯�S/��O�m��Wh�޽8`����Ӕ��V���֭���߯];w5ZOk�յkW�1B�ԳgOmݶM�4s�IR�~}�>�m����WJJJ�:�k�С��aÆ�k׮���Ү��ZUKbB��>�lI�i�2M.Y����Р��� @���K$IO>�wNZBC��c�ꭷ�Ҧ͛u�`��ٴ����=��|ٶ�[��	|CTj����{�v�_D�r��UOk�s4|�8}�U�����%�0�v�%))��Z~q�����	�  ��a����S^^���2߰Iz�W�_Ҧ͛e۶N4H�iʲ,EFF��+��[ZZ�U�V)55�o�����5l�0�]�V999��>UCk����j��Қ}������q�F�t�IZ�~����|u���Ƃ?!��  ��+���x����_�G���ڵ�BBB�n�:I��d�RSSu~F�^[�D��������w�ܜ\�޳G]�t�E�""�u˭�)%%E��ْ����_���˷�5�^��.]��q��N���}�Exx�n��V%''ש�5Ǎc#�� 8����zã��hM�:U۶oӦM��r���N;M�_v�o�����z����w��]:�
�$    IDATx0K���5j�&�_g��=�u������L�T�^�t��W��G�0~��9����Ou��!:tHOlվڢ�:;�Bz�2�[��ƿ�ܞoUQ^Ƨ �^����̙3����{���z5���_�L������	�a�r:I2����e�  #�@����ju    1F  W}��z�   �:    �:   @P   @P   �    �    A    A    A    �    �   u    ��I  <,�ҢE�$I�]S5m�4IRIq��x�Mٶ�޽{kܸq�Z׫�.���w���ӕ��ԩ���n�_�^{��Uyy����ԣG>B!!�o��}j~�j;v������a����sv���_�N�EEr���cb4r����� @Ӳ��UXX���m۾]�m����r�0�P���S|\��z�I�""":���?�HYY�JLLT߾}����m۶����:��3e�q�>~�9���			��ϕ���'����0�ٶ���GTRZt�� B���<m߾MÇ��;��¢��3�!���v}��	�>lx@j���UVV�"""t�g��phȐ!z������Y��-�m����:�III�<��tIҐ���pm�u  ����P�^��k�N��Ĩ��RCN���^sܷ��Ç%I]�$�B�i�JM���:�w�Ӄz��m[.�=�9s����^���XEG�(;;G�������ս{w4HNgpEc�:  Aj�����o�f�%��(.�a�1|�4F5�����s�p謳�kǎ:�uP�r)//O��0~<A  4-&&F]�uU��,�ߟ����(I:t(W�G�C�e)+;K����	��䅡/uTg������Po�����Z	�  ��G(�k��{�Tvv")99Y]��*++[��_]Ӻ);+[EE�JJJR���h� e۶֭_�{���U]�v�L+E�E���eJ��]����?|�{�OP  ͗���L��8q�֯_�={�j��-
Ӏ4|��N��-��M~�;;�G�G(�Gw�=��{���p(�G�F�tme�¹����r{�UEy�: ��Rff�fΜIC �a�r:�{���+-$�L
   %�:   @P   @P   �    �    A    A    �    �    �   u    u   ��   ��   �   �   �   �:    �:   ��	  ���JmذA�2LCI��2d��$���ڹs�,�VLt���[�Q�X�Z%%%����h�t�I
�$jÆr�݊��҈���z6mڬ��l���kڴi
���l۶m���TRR���t�u�]����$=������O������|Cqqq��ȑ#z�����-r8=j��ͻ��v�ȑ#Z�r�\.�bcb4n�x���I��/_���BIR||�N9�EDD��j_~���mۦٳg�Y�� l�Vzz��N��ɓ&��vk�Ν����2m޼EcƌѤ��;vtxMC���)S4u����j�֭�e7nT���5y�d���h۶m��[��7n\���������/ӫ�k@�Z�`�oٴ�����O)���ps�m[�7KK�,��E�T\R��_y����b�*:T�f�R|B�6l��[vꩧ*##CJHHк�kZ�$��䨲�R3x�1A � ����!�4������rIRqq����|=��]�u�����:dڶ-۶}�������\������={*+++`�HRBBB���8p@9���8q�$)#�<-_�·|��aJJJ
�z5a�9���hĈ�����z���UZV�=zH����={���GFF6�Y��ǣ�k�jԨQA�{��/  ˲�o�~0@����b���(**JYYUQ^.۶eF������*��WDD�N>�dIRyy�߰���pU�\�,Kf�F�WO ���(%9������*,,�����!@m����R�ogꪫ~١����*��P���(UVV�}G�/_���<EEEiڴi�g���0��"� p�m[�֭Sr�.JII��N:I��o�d+�*�utH���'�,۶��[��w�4hР�%F@ڧ�z:�s�a����z<����{4����0aB��D=ӦM�eYZ�n��l٢#F����<h�ȑA����/  SH_�^���uhjj�ƍ;U�ƍS\\�"��:�.�0����7�&<<\��e�����
	�����	���Tegg��mdgg+66. ��ͩǲ,�s�JH�ׯ����뉌��]�+I%%%
��1MS����w�}�zrsr�����_]����<��w�yGu  �q�F9LSC������T�w�¶��ջW����r���m�ڷ�b��}�'<<\��ْ�={�(�k׀�iiiJIN�G},IZ��?�:eJP�c۶x�A���jލ7vJ=��ъ���޽{%I۷oWϞ=%I***�նk�N�����VFF�f͚�Y�f�a��1cF�����I��p�]�_[nϷ��qV ��Iff�fΜ���)((��� ��O�I��6l�$i�ڵ:r�$)=�����ס����k��_���B2���i���~�3�߰An�KQQ�>|X�N��T=�|�rrsUQ^���PE����1c:���nۦ��p����ԫw/�u睾�9�|}���:t(O����ׯ�}䑀Գy�f�򪫕��$��~�F��;��}��S=bee�bcc5�j:���R}��G*��X:))I�G��]`���Զx�"����i'��G��$�p���9A �`	� �O�u��    A��   �   �   �:    �:   @P   @P   �    �    �    A    A    �    �   u    u    u   ��   ��   �   �   �:    �:    �:   @P   @P   ��4  �a۶m���TRR���t�u�]����$��KTR\"���c��;4r�Ȁ�S^^��\�~����.�@�^zI@������W_�[���\]SS����}�/_��_xA��~;WC�	X=���^z�%�=���W��v�""":�����J���Sii�fϞ���0߲#G�h�ʕr�\���Ѹ����wv=�-$z� >�����2��x����-��g�t�-]���CzS���oO��rk�״t�M�65`��$'��e�%�4qb@�q�ݺ����������.�P�?�D��9���'��y�a-��+�ѽ����^OϞ=5}�t9�u���X�JC�լY����6��Ɩ� 8�8p@9���8q�$)#�<-_�"(�)++�[o�����BBBd����҂�}�����Giƌ�Ƕm����r_{uI��zv��z��TJJ�$��q�lٲ�%''��k_\\�Ҳ2���C�Կ�ٳ'`�4�,�� @���QJr�Ð$������@.�K!!!��믿^�-�{����ZEFF�����+>.N/���֬Y���X��k5`�����$}��:a�`_(T=w�y���կ)�4�����z����{vkϞ=JOO���˕�{H�e�4;�϶��T�5BqTT�*++VO0�5  �mKU!�>ϟ�-\��[�B���'V���QvN������3t�m��}������g����r����/��zBK������g���{VOJJ�n��f���u���(!>^�����	�  �%RSS����\������-NKK�a���RF�y��oVOuou�8�I�&)//Ok��׶nݦɓ'��ڴi�*�+4p�@I��3�Ժu��r��>�&M��O�]O?���������H��������(44��t�:  �)--M)���裏%IK��GS�L��*���+��[��;�j@��'!!A#G���WK����k���+666 �T��|GS�L�;�'55E�о}�%I�~���{��;����ٿ�[K~~��]�@^xA�����ъ���޽{%I۷oWϞ=�%P�� �eo�k�k���V�e�$ �{)33S3;a(�$mݶM���>�W�^���;���l���M***�i1r��Ιӡ���z$iϞ=����UXP���(�vn�O?�X=�t���o�MC���%Io�����υU�4J7��|B���λ�n�zI�M/���;�G}���ڿ�������8M���+L�􌕕������N����z[����#�t�dT=���� @�u ǟƂ:C_   � DP   �    �    A    A    �    �   u    u    u   ��   ��   �   �   ��$��    ����?�/��  ZI���N���uk�!��
<*��.����94 ١��N����P�ߓ�^�  ��G,-\]���T�?��I�enm�r�
1t���dL�z$0�ߣ�Nh  �Vᶵ��r�{m�<V��[����J��ɥF����
u2�߳�^_h'� ���;�(��<O���l-��B�x�s#�E�:������   �i[�G�ZT��^Ӧ�n]��X;yh`|��z��  ���4oI����?e�Y��?%:\b����u  ��R�u�[%�k����[�
7ݍ �  4˳��kGn�Mٚ��?WW�� �  4e�K�^�y�y����A  �)W��x
ƶ(��^XE�:�   *��>��������B���?���&   8<������O������|Cqqq��#G��Ԗo���ph��њ7�F����I�3g����#I�۷�n��&%''�j?��l���5�9=Vg�PJ�Ce��?��ܐ���$iL�0��u����4��2��r�K���{���KTR\"�����;4r�Ȁ}^���z����駟�a����t饗th=_}����ۧ��R͞=[aaa����R���{��<�"##5s�̀�#I{���ƍ%��36z��t���	�� $�M����~J��m�:�YZ�d�/Z��b���+�G�n��V-]�DK^{M�SO=������n�z���Ke5��8:JC���h�_7s�-mIz��g�t�-]���CzS���oO��rk�״t�M�6����ٳ��O�.�ӿ_822R�G�=Գgπ�cY�V�\�I�&���֠A����_��z� Ç�����DM�0�V�1B;w�X=�����;���6S��fބ���$I?SgY��~=-V^^��Ίk��w��H��O0}������o�����_���:�������vk�޽:��[�a��v�j���$� �����T�ۙ��_��9s�jӦM��M�?�X��s��mA�4�;Ήק������7���_/ۖƎ=Y�]{�"#���߯��8���+Z�f�bbc���Հ�ڻw�����6�d��Ə�e˖)$$D�!�qƙA����  ��G�w�={�X_{ =�����|[cǎտ�����i����������X�1I��!u�u4�������������sTXP��=�d@�7�998p�,xV���Э����]�v�O�>���,m��N?�t�w�y2�$}��gu  ��0qϽ�*!!^�����t��s�����X���5����z�J�����N����Ք��&�0������7�����I�K�4i����TPP��Nii��9����֑��'�ۣ��IR�^����+�
�<�}  �ٶ�|P����w�����P��JOO�eY��|[}��m��"C����כ�?\]��}�!C獈��|����L����e��f%(�У?��t�� Z\R���d�\.��λ�?p�L4r�}�z�Ə����Zqq񊍍��h�ΝJOO���h���*..VQQ�bbbt������4ߟmd���E�m�=ߪ��L  |effv��q��ϟ��>�\��)11Q���գ�<�͛7�W]���$��!I5r�����';;[��v����4|������綥�^X�-YMϾ��I��?Y��\���a���HS���ڬ�%��nN=yqt��ϼ�ݤ��"���#Gh�9��G�N?x������PQ�Q��ܹ2dH�ֳz�j�߿_eee���P|\��L=:�̛o��SN9���z�g=;v���͛%I��!=z����:����9��`Ԩ��u  �)��^V�76�.�������#�0�uƨ ����������EP  5��S!��߈ilo�:�   ��54mPh�����j���  А��	�����0���Cix�  �#��#;/8_8*Liqu  ��\1>\'v��1�C�9tٸ0u  ��u���H��4/����T���`�r�[լ�t�6u�9Q
u06u  �fK�2�PF����K?{DV�!Y��*���&�O�15��(��M�:  @���г��hx��3��CO�8Z}�0.u  �V��0���(]vjx�s�G��'32YfT�"�ϫw���KO��D+1�؃c�� ���0t��p�7,T/���{�*T��{���_���!�y�rr(����  ��L�0-Bל����Z�ϭ�(�»NT���P�d�F�;uJo'73A  �3x�`�i�Bh�   �   �   �:    �:   @P   @P   �    �    �    A    A    �    �   �3'M  @px�����ǟ(;'Go������|��{�}���Kr{<�ׯ�n��6EDDtX-G��<�-�n�����Q�5oލ
�$m۶M����JJ�������Kqq�������z��5�3g�\�ٻG�Էo?�r�MJNN�z��˵j�*>|X�a�kj�Ɯ|��N����_j۶m�={����V�[o����J�!I?~�RRR�;�u  �Ĵ�����O)�V�;���'��y�a-��+�ѽ����Z�m�:�YZ�d�/Z��b���+��>�����2��x�������.�4Uk ���n��%K���4p� =����F���WFF�f͚�J�K�7o�[������J9�Ή�M�s�Yg)##CA�	�  ��Ç)))��뻿�N=�{��é��iٲeZKbb�&L� �á���1B9�9��('7W'N�$ed���+V����.�4Uk �'55��=nO��Oxx��w�.�0d��RRRTZZ�[��x�v�Z�5�S>���	Vu  �\߾}�{�n�ٳG�mk�����=$˲:e�����|;S�'O���	MIN�HMMUaa�\.W@�	���	D��sΜ�:�Z�j�����N����h׮]�ѣ�����k���:�%�H�|�7�xC�W���2A �c\JJ�n��f���u���(!>^���5�w�={�XM�0A��WV�����H���Z��O<��̷5v�X��_�:�۶��g��k׮�޽�$)//O�ӧo�^��#I�'Oֹ瞫3f���Rk׮%� ��4i��~��z��4x�`���wxP�,K��{�����󽞚����lo`�������8�����@i��@�ڜ}:�N�{ιz�������5r�H��99����믿��_]��;Ｃ�����#I��ђ������_yyyA�sϬ/  ��߯�ݻ+??_�.X�/���C�>���Pͻ�F�eiiiJIN�G}�ɓ'i���h�)�'�'�6�ς�B(==]�e)3�m����U�V��p��O�{����u�����-Ҍ3:t֗��q�\r�\����eY���?���Av�
5����|���2~� ��2335s��N���������С<%&&�_��z��G$Iw�y�֭_/�{��e?�y���o޼Y���j%%%�4��5r�������۶�?ܧ��"���Kw�y����VOcm���4Ukgד����n�]���d��>Qs���Cg6����{��7�hjj�ƍWg�ŋ鼌���SZZ�?��7=cJJ�F�����N�����1H�Q���_�:  A��Q   �A    �    �   u    u   ��   ��  &C�    IDAT �   �   �   �:    �:   @P   @P   �    �    �    A    A    �    �   u    u    u   ��   ����ٻ�8�����{�n-������;ݝ�$de��Q���"�>:�t�7�q���\Ǚy� �"KBLHY���V�[mw���I�;[w'�tu��~����uϽu|�Թ犈����W���L���>��˼��%|>�~ի�ԧ>I( �L��o|�'�|
�ir��s�U�0%������k�͖M$��TWs��?�������w�@ ���>�ҥK��>?�{��^l�a��Fn��&��pNC��'hjn��q>7��i*++ؾ};�������峷~���hN�J�hkk�u�@�ٳf��� ���`pp�ΰ`����SQ�qhkk#�LbTWWc�Sߟm,�&��7귇�l%�L�VDDf��kײf͚��Ooo/[�l�5�y���[oe��|����_���q�7���hoog���SV�Ѿ��;�;wW_}���Ƕm.]����}7s�����/�K������>m��|���?�UUU|�{���ã>��BGG���x���ﺋ��.n��f ������^�\�w��=��_]N�k�.���)���Յ�TWW��p���,v������'$��>�m�L&),,����`0DEE�	y�	���}� c����"""����X�j>�˲8�����̆���������	˲0M3�!}����L&y��ǹ��K��>��a&�d2�^�SV�ݻvQW[GUU �9�y䑜?���`��pl'{{kk+�]]��� ���oᏏ>�Ӻd2�MQ��������0~���q����~"��a`�2v&/^4�EDD$Ϥ�i��n-��hii�������g�_���h��~���p��)��h�ӟX�dI6�NE},�⳷��G>�O`�&����LY}�ݴ���&jkk���HWW7���|8��?�	6o�̬ٳ��׿@gg'U�������q2��e�,���1Ӳ,�����8�ϩ����<��8��y�Z�u�<�8���8��X�jU����NN9�~��������{�MSV��~�v-o8C��T�L&ý?��o���7��ｚ��SV���*n��n��K\{�)-)�g�'$�~��`���q�Yg��?φO� O7�����Jaa!�HDA]DDD�s]�/|񋔖��я|${����/��.���������g����m�΅^0��y�R���r
 ����cÆ�d2�)k�.�����������%K�P[[{�z��~?���2~��􎎎�����E��9�M��k;cg��d2�|�)�M�h}�����}TUV��k�����H�<�;��e� ���'�,+--���N�g���u�(..!�NI}�Y��A.Z��`08��S]]EKk+{�� ��OQ;wnN��x���2R�X,�~�C����O<�Osss��ڵ�����ٳgSUY��������r���9�~�?;<�QTT4eϯ����ކa�T����f}9�5�˖-[����������{���3�����&n�җ��S)�O�v����p����7����˧�}����?��~ "�B���z�,Y<e����ϲa�F`���k��ޜ�&wttp�M7��Ӄi,Yr*������6f����~��0�~���VJJJrz̒�$m�m��K 8vz���v���m��G0�vn��'�L�{�.|~?���V


�5k�	y�9Ҭ/
�"""y�E���EDDDD�s�������QP�t="""""y�EDDDDDA]DDDDD&�5N]DDDD$��Ʃ������aP�<��"""""��A]�_DDDDD�0��������������L4�k������Hu�S�à."""""
�"""""2Ѡ�q�"""""y�5N]DDDD$�������(�������D��Ʃ������aP�8u�<�"""""��."""""��.""""��A]��EDDDD�0�������T�	DDD�C?�6m¶m

9m�J,���g�ehh��H�e˖
���>�l޼���&.��b�������3��0FF�\�����)���8l޲���N0��ͣ��qJ�L&���Og�9�C8bժU9�O*�����u�fϚ���```��n à���p8<e���裏��`0Ȭ�Y����g��=4FDD��x��Y�`���lݺ��۷sꩧ�|�r�{���m�ضm+V���� �����dNX��>�sN�?�L�>[�n�s]V�^�a$�)�O(�ի��6m�DAAA�����FyE9E�"��������hko���˲��麟��y��MI}2�����c�-�����顲�r�_�yf)��������$�I���������=�|_H�<��>��u�V�,Y��O��q��ia��Ř��a9�m�q���`Μ99�O&����E� ())a```L�u���~���'�N��#߆�?П��"""������P(D:��u�l��3�>K<#.��3Ϝ��l߾���ڜw�T�<�PQ^��E��4��>���;v젷�˲X�h�htJ����������d�[��߲,���<�`���455����`1U�	��i��4�@���l�Ώ�n��EDD�Ñ��>��3�<��[��k�N-Z4%�����x��i�W���`�6/��"[�nc��S��>��L&�F�,^����֭_��/���@KKs�Ι�G��y���P[[K("���ږ�~8�ߢ�����6 
#�y3�Ĝ�a�\
�B$���1'�I�u��o�0���K��P1����e``�?=�z�1\�婧�bppp��g����O]]�xl��g_o��Y� ���&�J�N����H&������i��,���^�L&����0��$��e�)Z%��鐮#��(Rļy�7o�P�}S4��~䰮�v�\+(( 
���@SS�55�P�o������BQ$2e�ihhࢋ.b�����1M�s�=�H�t��ضM2�F�;���-*���	�����=2�IOO+��aBG��>�--��Tgg:�uP����q�X��������Τ�\����lh>������1���]������a�ț\,�F�������	DDDf��kײf͚r_���lܴ	;���0�ʕ+$�I֯[G*�à���%K����U�=��ì^���L�x��y����dlJ��8uɒ���<��344ĦM�H�G�F��d	%%%Sz��q�/_Nii�	y<'�I���p�@p�t��x���^ |�����?��T���V���ȉ��'�5&
��-b��|߇��A}����.""
�""�ꇜ�qt19�8�����q�"""""'6���u��u�ϟM�ޑº�>u�)�L&��144��8�|~


(++#��DDDfdP��9|`ׅ�D�Noo/�]]x�������?�@?�������DDDf󐉜Çu9���8]]�cB�h]]���q5����L
�Ƅ���.r���KgW��vvu�8�MDDd�����8BX7���E�ĝ`�v���a5����L
��#2�����ʧ�j4���G·��.�G<םTyw��EDD$���	�("��J���ň�Oj��x�q())���@)""2����)\a]dj$	�:;I$G��c`����~B�0��ՄB!5���������ENǱ���&��1e�d��ݻ)�SYY���WC���L�����Y�
�T���2��q?��ã�?���s��Qﺈ��4bz���w�npęE����i$��mghjnfhpP�.""2m���2ܳ�Ք���N�
�"����0��-xH��:���044���A��o����0��.�c�t���<�Ď#�<�ֶVR�����ȴ����K
qϘ�W_	�ú�L��4�ك{�z���aO�͹.""2����-^Cޫ�0��.r�uuuc�xL�x�L���n�i���a�3���w]a]d���X_^ԥ���d2��"""2݂��R����p@a]�uww������z�EDD�mP��v^R�w������Q�d2�׌+C����i����#3�,�>S-'2I��}��5��XLGDDdZ����b�����A���$��e���upDDDfBP�"!���*�Ղ"�N�ql;/���6�LFIDDd&u`d(���jA�	N$�~��:H"""3&��Ȅ���}%�tJ�4������@$�l�����*�"��y^�GDf�0�?
�"ӈ�8�]?��A����u�<�d2I:��ﷰ�>�Th���s]2��m��P�00�c���.rB�z~�X;�Q��s�!�H�I��[j���M�@�$�Ȥ����cY�H䘷�1�"'�����|�]�D"A*�$�("3�X$����/����������d��~K"r���-����M�z�EDDrғ�$����"'��qzޛ�6��T���S��z�E�؂��ևo�N��ZCDD�8u���>5��CPJa>��-�9^o�>�0���0 ��0��b��.��������i�5����}�����M����d��4FDDDDd���6�^�t(��n'FπZHDDDDd�����k�l�V+�����LuP�=0vtbn���p�Ҡ>&�Fg?��[-&""""rB��q��c�zs�.�DF�&""""�c�l"���2��;q���EtId������_�~���?���J5�Ȍ�G�ݜq07��]<��@-(""r=�̳�����5k��j���9f��a��t��ann����"""""��?d*�HϺ�anmU�����lܸ���f<�c���TVTT�嗷������0�mc�&�%%,��Ȝ9s�lo�ƍ4�����=�n��4"y�'6H}�C�ENv��L&�m{��!�a``�2��O(�0H�<�a�v��	@0����֖�;�z{�H�Ӕ��b����1z�������TUU��P(Dgg'���|�Ӡ~@�@"7�4Ղ"���;��6u�dҴ���a�[TWW�Dt@E�X*�b��] TVVr�y���O���5����O#��dH�Ӹ��c�=F:�������*��dv{��՜s�9���O>Igg�\$?���º�4�00�Կ.rP��Ӳ���ܰ����̛7�`P3<�L��xo�kJ]]m�ۮ��ڃ�zG{;��lfxh���$�	 ���ۛ[;so�[m]���H�uoo:?8���a��<�=��E���kڇ��+�������9st`E��8�o���M���j�����y�4��������$S�Cv���7v��3�Y>��F�L�����a���2h�������ڟt*��*2Ţ�h6P��A?�7=�e{�O]����:�����c/T-.�n�e�<���<�����"yf��c$���`����nv0��[d���f�\����頊L�P(D}}=;w�d���$#CX:�%ť�|&�����^dV�,����c߬�� ��ر���v���wxx8����3�i��}&~ˇ��������CWQQd��O��HX�r%�X�EwO�i�|��1e
#��q�YD���������(,,<h{+V�d~c#�ea;�UU,9��Q��,B$����~Sv@����/�GƦ{{o��lhx��'����<ϣe�������2w�\M�('��kײf͚I��8�X�!9$�I|>�ee_��~�i�����L���7���u�E�A(�P�`(�߷��犒�����w�4/�Ǟ\jd�fU9蓯a0g�\b�8C���d��$RTD�q�"2�tvv�~�z��J�,�X<��)f���
�"��|p ?DV?촍z9TX/-)���D�!"y)�RZVJ<�O&����SUYICcØ+��H>�lX7�N�4n��馤��ο@!����A'�f�b4�&uə�y�\r���\2��G `v������G?��g��ZQDDd�������������B~�aj���	���C__�Q�_VVFee�RDDd:u��p\�L�����m�@��;^��KE�Ǵ��EDD�{Pw�L�ƶ���m��c��a]D����B8�{�<(�Ո"""Ӝ�H��ҳa=c3��Rԝ.�;ˢ�(/�)*:�yɃ�>т�a�%L�EN���*�I�j�>��*�x"""'SP��_?Ԕ�"r\f��`{��ɬ�,K��"""'aPw�b"'P$RDmm��۲���QTT�F�!��)�y���|��t����444000��@?�T
۱�������)*�`zF�����A��8٠��.rb�A4ZD4�s���9�<��v4FDDDD$��:��q�r"""""��]��u�EDD����u��r.����׿V����Ѯh���_-(""r}�;���~��?{[__��o����a�|������ڴi?��/��7�N}}=�@P@$��G���8���ɡ={��O�+����������)**bٲeD"먶��Ί�W��%��)""�3ۼ�[n��z������A�u]��~֮}���N*+���Mo�]�";U��>�y|>u���}�!���Y�l�_���|��x��?p�%��W��%e��<��C��W�fOs3e��:�����p8�ݶa̚5�?<�zz{����/��5�u�T/�_|����/��
��1���k�y/��rR1�ee��8u�\x������������|���~�s���}\�Ϗ�#�}��}����7���'�x��㞟���~�S�ַ��gn��O|����?<���e����o�|�.���]���?���/ۼ���y�m?�䓘���w������²�^�H��m��n��%�.�w}���|���D�����12���㭧��/|�6.���\���}��<x��\q��Y��9s�����Ov�x�;�ek��򞫮 �x�[��׿���ޯ��sϽ|�ൗ\��Y������е��/Fii	 UU���?��4'���588��� g�u�f����Z
QP������ȃ>�E�Ws�)�d�uww388Ȋ�Ǭ�r�J��z{{)++	�u�cʔ���H$H�R��8���F<�_��5��k_;hykkK6l7��gC�d�=R�JJJ�����o��NcŊ�:�\��u�Z�����n��/��u��;�t;+V� Fzԁ�X􃌺}t��pS,�$�+_�2g�y���z�����O�3�_�N�}�9֭_��w�����\y�������&�?���go��/��n�����W *++�D"lذqL�6P\\LYi�Q���ٳ�F�<��'t�Cihh��+.��w����z���W
9�G]DD$O���?��(,,��[o��o��.��ﾒ{﹗��j�/_���/��_��~��t>���^����ߥ8Z�E�Ʋ,���x��?s�7�d�њ����Cq�s�������7�P_��(����H�0��~��F�җ� 1��]W\��8�s�O��ꢪ��k��������|o{��(.)�W�����/���̙3�U瞓�u�	�C�nj�G�/�Gq��3�8�k���r>�Y4ɩ[�Q�=lg+�dB-)""3�ڵk���L��8�b1
Հ"'�P(4�r�P�o`��!�[c�EDDDD򐆾�䡁�Z[[��744TWu���N�ٹsG����R]�BDDDDA]d���|��ƶn�d�UDDDA]DN�����|*2�q��|Ӣ��c?EDD�eF;�x�d2I__/�t���B*+��1�z�Goo�x?;��(**�����;wb� ���̞5 ۶���!�N�Ngp\��0M��5�~ii)�1��'����.zzz 0}>�_0�j����ʎWpl���2�����=00@<#�J�8�a���	,� eee��c�މD��X�D����cw    IDAT��� �H!%%��?���$��bqR��@����#�u:������T��:s��� �d����l��<��֖1e3�4��=$��g3:��i}��:I�!�L�PWW;�^��n/-�u�q �f�ʆt����q����Ggg�A�6��d��F�n���ؒG*�$�J�ǩ��;�I���g�?�.��x��9�_~��&�������i��>��v.�[����V,�b��%446Lxy��a�/���F*�$3�|,X�W� ��.'���A,+@(bxx8Z3�4�G����cB�o������>,+@$!����<w�w�o$Х�I�������P�'��@�������! ������'4[Jo�� )�-*��f�!�L1846���	�E�(�����#�ώm�g�����6<<��oQX�4�q�y���~���p�%K����2������GII1~����6�J%�t��x�'�F��W���<W�0wn-.�
�/O=E4ZLUUU�새����B���u���mۼ���F.��Nd�[<ˮc�&������

�ho;��� ���cn�<����fp` ����	���^qqq6�b�6~��uǄ���	���9ٿK��F*�yި`�3&�Ϟ5{��iA;v��˃�����{�y�F��L>��c?E�Ŝ9s����Û�r�qx��Ǹ�K�F�475�j�y��̝[��&�+��<��s���_PX���gp`������u9镖�g������g������tj،D��(�F��h����```���8É����Q�O��h��a�������� �%��#�h�|���T��Ϟ=XV`��� �P�Ha�M]�%�Jf��g����H�R��֣������t8��c?E��M����/$�04<��8GGuDinn��:��\����Ʈ];I�32�v��u�т��'�H�z�ݽ'�cpңa��~�L��zl��;���A��(;vz��oP�g�E����դR#��a�'|��t�������%�&��m~�G(<)����O��b��#=�vf��e��Y+��0��\[�h����t���כ}�O�}QP���26�z��%5M�ad�ٶs�:�!zH=ϣ��7�8f֬���~à��������z,�+--��D"A"���Y^<�z$�I��L�t:�p"����tuu2w��'L�RVVv�m��q�e�Iq�՛.3�����0���L:�}]o��|��C�~饗]��~�~?sk��������Y�hQN�ADA]万y�@ ��1848fn�X<v�a�mg�� e_�=�3��D��� �P�drdZ[[�˂�����ql|>?�p�p8��������N ��T6t��l�QUUyP�<����	�9���t�.��lfႅ��������P���D��2����'���l�E.�Ad�QבLţ�-t�]�v���Ak[+]����=�^oo�x�������c�'��s,�+)-*3�ܷ�سg�v���X<��� �x?����b�o�g����=�L�ݻw��188@<����;w��ކ�:�"y�]��������Y�.���
�T
�0���c�K/��d���eO������<W�`�6/��2CCC��iZZ��{w��y�"�@=�2-�3<4�=�Ҷ3���B���N��/��AYiYv���оw���#�H$&��s�ۋ���1���0����yd�??\=�������(�L*;�{:����]�[$Omٲ��[�f�ߵs�,:�eK������󖷼%�lŊ�<�n����,�eK���e����0���ॗ^±m

Y�l�u�����"
�"�ɳgϡ���X,����}���r������lY�o�E�����z�HgҘ�I8�������I�cٞa�D������,�Mz,eyy9CCC$�Il�Ξ4���	PZR2fH@EE%�H}}1�al�ή���(((��0������bK�.e�ҥG�|̛����g�u��s�>��s�]5�2E� ��,�&��7귇�l%�ԛ��뺇<�opp`�E5f͚=�B��-r,֮]˚5k&���Urc�ENR����?���}���8�=��Q5�L{�����D
�^0�a�f��wK�����e�dh��<�<�-��s�b��J�[DDDA]�D)))����J&q�^�4M�� EE��K4��������ȉ��j��������A�Q"""""
�"""""��.""""��."""""
�"""""
�"""""��.""""��."""""
�"""""��.""""��."""""
�"""""
�"""2����|�-��&"3�_M ""�?��������A�_vٛX�t)�dB�$��."""S�����|��cn+..���B�#��."""S����3���n��ί�ǹ������>�y|>�,<����7���s�ԧ>�3�<Ï|7���,]��o����r5���������=�<���۾HOo/w��e>��ϑJ���'��0M��/_�[��6�����`"
�"""2�]]\|�k��v�}?����H�O��1M���%_������_���� ��w��w5�������Lԡƨ���Mx��c��'v������"��ݖH$H�R�A5����������|�1�^��ۻe���� �u]5�H��<�"""""
�"""""��.""""2M��ɭ���a;[I�*i""2C�]��5k�Lj�q��b�ENR�PhB傡0~�"���C��z�EDDDD򐂺������������(������(���������������W�����uٴq#�$	"EQ����ٳfe�ضͺu�ikkŲ,�,^BCc�!�7^��l�x��D�q��ADA]DDD
�g�}6�p���V������߽.;'��MI��\�f��<�ԓD�Q�+�q]���>JJ����G,;޶r�Y>�� �/4�EDD$O��~V�\III	�`���
���� �<��f�,9�` @yE9s�ֲ��	����?���иe�[��}oy>새�����Q2�d81L�����aǡ�8�-S\��?��^x!�Hdܲ�-��>��<�Ad�>��	DDD��z<��4�7PTT����,+[�
X8��a���O��x�s��-Ϸ}QP�,��x晧�AV�\��M�y��d2�p�Ig��|���Sv2�x��y���^:�}���\새�����5�uy��g�<8��31#���� ��G��9�'-ή�y�f.X8n��O4�Ov�[��}�n4F]DD$Ox��s�=O*���3���<\���<`dXHmm[^z�L&C__-{Z�WW�����
�Tjܲ�-��>��<�A$_��I>G�������	�����Hk׮e͚5�Z�qb�XvJŉ���:��+��`�B`d���׭���mB���d�u��a"�8�� r<�B�	����}� c���
�"""y�EDA}tP���<��.""""��."""""
�"""""
�"""""��.""""2��ʤ"""92r�M���]�GD��s����գ.""�#��DDA]DD$�dlG� "
�"""�&�J�DDA]DD$_��a��C*�T���lғ��C�����H�z0���H&�d�j��D&�f81��.""��A=
��� VϺ�I �L188t�f���"""9
�e�8��0�H�L�	�,?��/"ӛ�8�36�T
�u0#�!]A]DD$��I8 ��d{2�@��"3������aY�����H>��|�y�d�T*����P��M	�B�"""2����`��au����/
�"""'�M\Dd���"""""
�"""""��.""""��."""""
�"""""
�"""""��.""""��."""""
�"""""2]�TDD��</�#"3Ͼ��++������x�G2�$�N��[X~�i*��̀p�.���m�P(�a��\QP��qH$d�i��EAA�Ed��u�$0	,2�4���X�E$9�mk����H��K"� �Lj��
,���qٞz�EDDr��<2�V ��o�ADN~�E0��m�G]DD$!=�L�y�`P"r�	�罂���H�z*�RO��(�����[P�<��Sc������H޽���6+"GO'�������4�+]d�>�s���G}�<��.""""��."""""
�"""""
�"""""��.""""2�izF�i�������+W�a�.��B**��]���������RV_t�a˵���ק����ϧ��rBu���'Z�h�z�"
�"""3�O>IgG>��o|#�e�Y�ק�JKk�i�f��� ��EMM��� ���XjLu9^������q]�����ؘ]�J�iko`VM�`�h4ʹ瞛-WSS3��x�����l���ijT�(�����8�g�&�L�hڽkLPonڍ뎄�y�� ���v���ƶmLӤ�����3g.0v�GCc/m��pb��/���up]��7��܌�y̞3�ʊ���uw��e�f��8��!`(*�2�fϚu�m����ho���s�8Dg玝�޽�x<@���y��?�ad�555�k�Nb�8��P__ϢE�&]����ڴ��XdQP�iàv^۷m��/F,��d$����@8����ޞ>R�4%��X>?�x���nz��9� UUU�m��q�~�P�!5�mظ��;v�ho���uL۶y��'p���b"��'�v�PQ^~Ƞ�.��_��� �j�*JKK[��6��+/
�0M�x<�ƍ����q� ���ٶu >����(���t����p!�0���}N�ME�EDDf���F�o۾7�d%�X�x<@}��l����O#��dH�Ӹ��c�=F:����yLPw\��O;��Ɔ�{I�R�ڹ���J�;�< �x�	����円�p�3�8#ۋ�.�T��:��S���B!�;�<���a�`xh�Wv�@MM5�y�9��ɳ�=KsS3MMM,X��`�ʶUiI	��;�@ ��y��㓪�D�s�����������),������.���X�|9�v��p�A}}C�lG{;��lfxh���$��1��B!��9��x<8��j���jk����"


���e�F���d��m7�C<��4������b}�z̝[��]7��榑o�z{	�r�����WR\2�zL�>G����ȱ�"""y����L&CsS��{����p8��� �?�<�CÔWTp�gp��g�{�����p(4���^�0�G�$M�d���,^����j� ===���%����m���#=�[�n=�v�&pˑM=�tiSu�d�ܹ���7��d ��W�-�Ų=��.^L]]���d��!�9��h4�-7�}�� ���86��z*�Z��_�z���������[��b�
 v���/�?b=JK��]߳��uh�Ӽ�LYe�e���ܱ�t:=�=/{2�D�1���l��}�3�i0����/��m���0�Y��^,).��3q���"�zf�Լ';3���B��׳s�Nv��M212|�󀠞J&y衇�D"D"���IWW�H�J���`�6�7ofǎ��L�����`�^~�e��;x��1M���!>uuu�!(OYȶ�����c�ڵD"E$Ô���jԴ���c2�)r�^�"""�g������3Gwa��3�<�h����~���X�pA��GGk�ʕ446`Y�==�����Ɣ�j�j���^:::����ϛ�k�>���^�x1��a����lzq�aˮX���O?�Ғ2�4�d���bV,_��_��l�eK�q�gP^Q�a�cY�哮�D�S�D1M�7귇�l%u�	+"""3�ڵkY�fͤ�q�X,v̡YD����a���}� c����Q�C
�"""""
�"""""��.""""��."""""
�"""""
�"""""��.""""��."""""
�"""""��.""""��."""""
�"""r��y�W���[�"S̯&��T����G��(���afϞ�9��{�����w|��D�/~��cn_�t)�dB�$��+�pϽ���˯�����e���7�1��/~�K���q�m|��͗]���0_������x��^7���ٰa����l���m3����������y;<��S���g��,��F�MA]DD�$����+�<�,��C�r�)�Riv��ɶm�NX���7�@��v75��O2k�,�� �t�����򏍒>�@&��g�����Lx=����Wn��3��K(�����۷�;�JwO�����8��ә7o޾O�1QP�����?��������K/�޾d�b���5���{�y~v�}�ڵ�t:ͼyu\s�5�u��2������|��ֲ���f��e\�u����/_��� .����^�;��*�x��o�m��g�6߿�.~��GH�R�}�Y�\���������u]��~֮}���N*+���Mo�]��0� �bg�y&��_�����k��>����X~Ŋ|�_�6��o��~������ٳ��w����n��f�y�Y��^���7PRR�Ӷ0MӜ��
�"""y�0**+ظq#���� �]�&�ϟ�i�<�����[��]��O<�W]u���'��)n��f���o���}�O}�dҙC}9����O�C=�u���/�/O?��w�d�v��Ϲ�g���+V�`�����7,��;��= �X$�T���l�o����ܹsx�e��׽�4�F�����@ 8��ZZZhn����&[�K.��g�y�t&ú�����r��7of����x�b***�EDDNv7�p_��Wx�;�Icc#K/�3^͹瞛��[���1�\}�լ_��>�'�����k��fǵo~˛��׿1�:�w����_�����lٷ���lۺ-�k�y<�s���
֬�v`Μ9����ӟݧ�>����K/m套���+��я~�0���^GGG�\iYY�����ߣ��Bcc#�p��GKK+O<�g.���Ѩ������l�ҥ����+��͛�����v��,^��;３@������￟��^$�a;6��TWW��Vm]���JKI$�R)�����4��uuu�H$X�l��N=��lP���fpp�+��)�r�J��z{{)�$�s�9\x�������u�]OWw7�����}�{G����/���u�����;Y��z *�*9��󩩩�._�h��=���(��������`����7�7����:���Gy��^�M7�LAA!�?����@0ȝw�I�Ό����غ�;��L��8`���wP�:�Xt�Q�6jk����ټ�U�⡇�q���)-)��w�����w_�{��jB��������ۛ����;���H�ECc�G,c&��MI[ku�<7{����c``�m۶s�{�b�ʕ���PR\��;>��q�Xf"�WYYI8��M/�Yw��-c�D"6l�8�̆(..���Tz���{رcG����V֭[�����H&�$�I2�̄כ3gN6����288���� `Y����s�o�����L2�$�N�k�N�;ڳ��M=�"""y�C�~��^r	.������N���}X��ל�
)--��<�ʕ+q]����tvv�x�I X�n=���().&. �Ɣ��������|'��?555,Zt
y�i�����t�0x�����{���˗�~���W����|شiw~����q�[�n�=W_������y𡇹�'�PPP@II	����oi�uŻ��8�Â (+�4�� >�p�ͷ����ﺒP(D,�=�{wUy��3������EP�.���
��VA����z�تŶ�h�Rm�U�]k+ֲ�"��HY���>�?C"[�$���3���9�L�;O����:�K0�`w_o��@ @LL�9�ܰ�2��.""�	���_|�o�A}}=�q�d�҄�    IDAT����'3#�x���~�)S�b�;;6��.����t�Ulٲ�ٳ櫓���
�mY�-��LcS#�=�8�����M7�Ȃ�Ce�M����g�)//�w��̜9�뮻N>�\n��+n������98���[nfŊ����SQ^N||��\s�drrr��d��ܳ��Ֆ� �=�G��_!//�Ɔ�u�^�j�Ұc���19sL����&��1�Ͽ��^&""]��ŋC�����罹�����n��|��l��ʳ���D�n�n�������lʦ��J���h~T���������b6o�̈#0|�z5���}~z�O�sDN�������2���{��O��)�� i���}�]a� ��."""r}���?�Y;B�ixFuQPQPuuQPQPuQP���{�9s�׎���"""���v���o��g+�[T��j%55��F����'::�M�9��3q���C�M��߬\����Bj��qFE�����'�_ܪ�ƍY�������������k���.�����̝������Ky�ͷx��玺����'Mj������~�JJ��X,<����*����tw������{ؿ?7�x#C�&::���B/^���d��)mZ֕W^q�@b6+
H�w-b�Ν8z%$PRRBMM[����j�L��/W����E �n�㌊bǎ�a�#TTVr������e͚� 8��z�o�w&�)��-�?U��~pĴM�7�v��|�D�����U����+������Hw��_��ޢ"�������^�߿?�q����� ��W�x��W),,��񐙙�̙3}y��{���Z~�ۇx�0��Ӈ�>��ʪ*������&^}�5/^By�~{3骫�6m*�A������뮟1d�`6l��_��~
����'���³���trߜ9�Y���r�W��>|8���ǜޖ���ŝR]=>��׃� E{����Y��z�����={�EDD�3���G}�e�]�*��t(����3i�U������'�|̜9���_�Bff�1ױj�*�N�ʋ/� ��b��_��W^�?���Ç�a��<��SX,f���z�n��[om��aðZ,x�^��� طoEE{���a]|�ŬY�����?n���' V���r�rs��I�L&��R�<i�^z)F���˟0~|X�ACc#~���ؘ�k��1��c��.""!���q�\m�;n��V?Ϙ1���O>e��[�9_��I�v�,����$�� ���S�Ne�ĉ ���RRZ�˯���ލ���[x�^�F#7�t# eee���={��'�:��\VV��`8��('����R�򶑗��]�v1{��6/�d�Y����� ��~)((���.����k	�g�Z��+����t_�`��e���x��شy�55��>�ԓ��t���fe�B:@EE���>�U�#F��k�SUUE��I�>���3����E�0�M�{｡.U-Oі�k p�s����g�؜�9Z\\��w���
���"f͚uJ�?�g�$h�����}~����G�l1�������x1�L
�"""�Ybb"v�������o���(��ɏIJJ�j�1o�<�>�q�ڬG�rp�>��ޭTTT��C�uk.={����Ͱa���%'�"X]Uz^YYz���D]]7��|��M7���[n!==�պRRR5jK�-���S^Q���[�s��E���U�(���D]]������{Z���Q���	Ƴd����w�25558p���w0c�-�1���d�bcC}{��� ::��7�z}�ƍ����3>^��ظq#?��Oغ5����yv��V!��E
�_|����z� }�q�A��Q#Gq�\�\.���/�, ???����b֯_08�蝘��凋�` ==�ܼ<�^/����ۻ�̌��rLԢ.""A~t���n���wrӍ7r�C���
�x����p����Ǳz�F�A ��������3xpv���M7���INNbذal��5�����?��F�	���عs'��2=4-�G4o�� w�qs��Oqq1S�݈�n�F4}�t��⨯�g���{�j�:�d�2^|iN����8JKK	 L�:-Ժݖ�����X�~=�����X,=s�i�EA]DD$���у��~���~��>���^z	��Fjj
Ə��+��h4������0e�T�vc��p�E��:�M����g�)//�w��̜9�뮻N�	r����_@���Ru���<��<��
yyy4640`� ���.����`�_�{����r3+V�$??���r���HO����'���Ӯ埪��c�5�͜7ztD���`{��� >�6ܺ뙈�tQ�/���V~�����Аv"�����6����Mـ��?B��.""""��EDDDD�EDDDDDA]DDDDDA]DDDDD�EDDDD�EDDDDDA]DDDDDA]DDDDD�EDDDDDA]DDDDDA]DDDDD�EDD|�!�>��v�Hc�.�O?�4+V����_��������Ʀ&���!�n`�ƍ,|�ers���|dfeqݵ�p�e����ڵ��s�.JJJ 6t(O<�x�Lcc#��;�	��s饗��o��s�u�w��3&O�Ԯ���?���������I-�MA]DDDN+�χ٬�Н|�z5���+� v�gT;v����������} v���ʕ��ӧ6���sĲ�^/k֬`��A��,�:�LFS���T���8`�Q��9����C[|ڎ�ށ"""쫯��ʫ�RXX���!33��3g2��s�9Oii)���_���ɜ��iӦ.����`0ЧO>��#*�����K����p� �[>Of�$�͟?�@ @JJ
�����}s�f�Z.XȕW\A\\��=�E�����(fΚŞ=E�Z����y�O<��8���w��F�����WP�`���L�t����h0��'3g��<�׿�h�;l����7g�Ǎ�'?�	F����X�jS�L��_ �n����������%�m߾}����Gtt4 _|1k֬����~�&��v<111,z�� X��V��rs��I�L&��R�<i�^z)F��]�N[�ne�֭��у�������."""��7���3f�`Æ���O�9��VӾ\���sf歷2e��^F��I�v۬6�$�g�$򕕕�����z�Ы�Q˜��`8f�wF9q8����������m�ڵ�ٳgw�v��f�j������!��� ��/� �~��aw�1�L��W�ʕ+�0�bbbb�EDD䰪�*^{�56m�BmM>����$%%�*�e��/�����\z�'���YYm�s[�)�C0�����`������g�؜�9R\\��w���
���"f͚��q�H? ����}~��t��|rrr�yvv6UU��ۧ�."""��7gNgw���$%%a�٘7o^��U���tz������3f���˰ڬ�]�9$'��U]Uz^YYzޞ/auuu�xS�E�7�t#�o�����VeRRR5jK�-���S^Q���ђ���}�B��c1����r\4����H�:p� ۷�`��[1b�����Ɔ��˟��G����o���۽��1�M����.�RSSCA��/WS__O ࣏?n�g�0j��6//�r�p�\x=�_�,X@~~~�Lqq1�ׯ?�M�NL���h/��Oў"\.��J�JIIIQP�â�����c��5�A�~?}�y�����111���G1`��_�Kmmm���m)))���g��=�����xOy�����F#���L�v#7L��ڵ_0}���H+�7of��L�1���b �m�z�����Ā0` ={5�5_�t?���\5i2�L���[gR^��R>m�P�v[�#�� ����X�x1��s�a]��니�H	����F��x���~�)S�b�;;6��.���~޼?p��~��~�<2���hi�UW�e�fϾ���������L�L�ͣ��c�˯���GcC�k����/�s����W�j^��z����_�{�U���̊+��ϧ�����8��3�������{;NEvv�у��LΘ��9&���tl���߆�դ�[DD��ŋ3q��v�������!**���{�������O>��/҉���6����M�4�X��͕���EDD$�ݻ�%K����՜�����"""}�3q�D�M��""
�"""�����N�V��EDDDDDA]DDDDD�EDDDD�EDDDD���bR�01���G
��I"��=n��բ.""&@;AD�EDD"����Nu�H�v��DDA]DD$R���˥"�ݾ��:�K�����H���f�d2��r��z�SD�	��CcS�����H�u�ݎ�d���Q-�"݀�妾���F����"""a
���ߏ�隣�	�ۃ�f�j1c<�E�s��x�>�n7��������.""��F#� ��
�.Wj\��f3&�	�Ţ�.""�L&N��`0�����v�&G"]ԡkS�v������tFc��`N��á�.҅���EA]DD�;�i�}�uQPQPuuQPQPu9ݙTDD�;C�D��9t�Ꮌ�����H�� .��ǃ�l�b6a0�E�@8x}~|>V��ݎ�`�h<��+
�"""a���ijj���`�Xp:��)"]-��X�F�V^����:,��ѧ�l�Q	�@ @SSn��͊�j�N��,V+V����!�S����H�A�^/��٢"�M��l�@�,K-�"""a�.��`0��f��f���WP	CPw��jIu�H��`�٤�!"
�"""�!k�Ǭ��<]L*""&�äk�t�����[_�EDDDD"���������������(������(�������������H��EDD:���J>�l9#F� `�ƍ��%!��1��W\��/�`̘1$&&jGJ���u�=n.���S^�W_}E]]-&\�G}D\lg�s�����Hw�r�*���a2���+�X,����r5���a4�8q"6���Brr2QQQ $''c�Z�3%"m޴�;wҫgOƎ�jZCCK�.`�����ǟ�m�����q0h� �v�i�_
�"""�oV�����)*��~�in����b �$'c�� ���iՊ�����ow0$b4�G����f������Z��bC����t:ill<�ۗػw�yzz�i�u������f��v�gwa��^�g7�@�]3�� عsEEE444���0����1�?RS� lڴ���"�� )�)$&$u��w裂����Z������g+�?��ʊ
z��ӷ__�r����Ȅ	����A��O���II�s�Y#C��ݻ�?` [��ڪ|Yi)�w��@ @lL���$��s�u�Y����رs^����F�Eii)[�n�����^�8��sB���`��۷SPX���	��A߾�4h�����Hwf0H��`��TW״jqܽ� ��ARR U�ո=��㱘����PYQAeE]d�w��lܴ��� l6+e���+>bݛ7ofǎ $$&`�@yy9U_���v3`��V�kkkY�n=v���.:"'�7�/�>_�С�0���+�h4���|DP��|���K�X{���r�j&L�@LL�1�QVV��h�/���b�ڵ�^�%�@��G��`4�n�z6m�����`������qֈ�JL��l?�6m�h40`�@u�n`��c���y!qq#���������L #F���j�����x,_���Cў"bcc),( 11��.���+WR^^ZgSc#;w�`��!9c �6ob玝|������d
��y�H���K0ԁ�v���3��=E��ח����fa<xn��������C�P^Q�޽{9�3����¨�G5�_b!#=������Pױ��i���<۷og�����ZE��KCSyy��EDD���({'R���={�0l�0
�[�YY}Ce�JKٚ��Ɔ#��6������茌�P��HOoԫ��C�r�r���m�,��O݁��Ņ^������7�]"핕���݅�NJ����s�=��}D9��Ͷ�mTVU���`�׋�u����Ʒ:7�v�=��6;>��ߏ�����1
RB�^l߶���j^u��`2�(�_���h���������� ����u��镐@߬,L&����M� -۹��z����pɴ�T��G ����g�i	C����L�ٲ��&99	��~Ԡ���UX,���a�d2�n�z���q�o8��ͦo�v0��A8�_�N�_�ty���H�IMK�z0oܴ	��@FfV�LMMM(8�1x0�����*jQlق��9@||�P9����3���e�&�G,N��[�F��rj,ii��߿��_�Z�x<T��0x�z��f��@]�o����b�������j���aբ.""a�F��ع��4w5��b�Ÿ�xL&#~�-�l�Oe���sh���,


ؽ{7��& �+�8�N����Ν;ٽ{7��5DGE���Hm]-N����/"e䨑6��z�0o�Y))-!!!�@ �7[����E8�Y��Mn^.QQNz%4_L�k�N�z�i�?
�"""(3+�/���n-�)����sG��5���:�/bǎ��ׇʍ1��h/��$&&2l��V�>�ؘ

��������y���>): �/��c�th�����;�M�7�����d6���J���x*H� ��y�\_�p�r���B������7��A|�m�]M:�DD�KZ�x1'Nl�<~�������BE��ikW�݁ٔ�#��>�"""""HA]DDDDDA]DDDDD�EDDDD�EDDDDDA]DDDDDA]DDDDD�EDDDD�EDDDDDA]DDDDD�EDDDD�EDDDDDA]DDDDDA]DDDDD�EDDDD�EDDDDDA]DDDDD�EDDDD:�v���H��z�̟�,k֮������tn�5���??T�w�a��ep����������&�����/�����7�ɓ&�yz8�Ж:Fz �|��|���TW�+!�k���)Sn��:t�z#���~PP�"|>��_��~{�r�Jz�7��oϓ��
@BB�͚�'�|z��~��-[�0h� �̟OMM-���
EEE��/�oVÆ8��p��D�;C ƏǴiSq:���˯�k����9�uh�r�7���!���B]_DDD"����?��A�ǤIW���Ď;Cerrr����GTT��755q������G}��[gǰa�?~K�-���MWN4�3�`ذa$%%ѣGR����t��x_���T�����
�"""]TUu5%%%��׷M�N'O>�8�������r��߿hz���ٽ{7�	�Wu����T�����p7L���``lNN���T������/"""�����ÿ�+�"3#�M��F�
4�&Bs��!�QQ464�i�wQ��M�Lu����s�Փټe۶m�錊�:��z;C:����Ԣ.""�|>s��%..�;�}R�88����Q�6Mw�R�H���� 11�	���v�y�7#���H�Cgz?(����t~���?L0�_��������>�<UUU$%%a�����M���'33����Y��M�,u�� AJJJ"�����P���~PP�� ���﩯o����� ��@ �*@z-��x��� x���R[[��lf��X�p!`kn.�|�)�]z)�	���'�������;�Cii)��>�e0r�Ȉ�é��3ԡ3�N��@v�}�[<����v5�7���tI�/f�ĉ����SSSs�Q(N��������Ͼ�'\�� �����˯��j�M7����#�k9.ttt4�L���Fm��8Q�R�H�������"/o��&RRR�4�*���ڣ.�tԡ���u�����no1��  �IDATS9�݁ٔ�#���.""AA]D������"""""��EDDDD�EDDDDDA]DDDDDA]DDDDD�EDDDD�EDDDDDA]DDDDDA]DDDDD�EDDDDDA]DDDDDA]DDDDD�EDDDD�EDDDDDA]DDDD�;3k���tN|��Ǭ[�����Htt4����:�,��4��|�\���+W���GUe%���I�8` ^x!]t!f�Y�Au8!���`�f	�x��o��j�oK�/^�ĉ�5��罹�������W_{�w�]DCCC�i������"Tu�:|�ʕ+yf������\jj*?����3Fǡ��n�������l��zT����H'���_��GYY�Q�B���wi�����o���}���2m�T~t���KG��.""�I��_�����Yf�y�U��-��ƛ~t��::��J����t�����;n(?n�������O*����o�r�J�K
�"""�QnnO<�$���/+KJJb��l��;x���Ny9�}�ϧ�ЍϥcQ���r����~צ ׿_?�!Ljjjx������-*�l�KQ��S^vqq1+W�bܸ�:ݠ
�"""]Ļ�.b߾}m*����:����.�G����eb������?�<�A]璂����t�������-f�������sO���Tm߱]ǡԡ��G]DD$B�[��m.��1�U�SSSS�#�>��P^^���ꠠ.""�E�]�U�ʗ�߯:t�w��G��.a�������_�^��Ѕ렠.""�Elڼ�]�o�����v�:|�����6l��}����W^�q�uPP�"*++�U����M�6���-v�`0�����_�^ǡ�AA]DD������յ{��˖��`8}�����t�X�EDD��`0x».�|HYY���RSSOj��Æq�/~��/�d�Y�d	/��"?�яHNNn�2rssu�XN��g��h�����v�\ѣGfͼ���ա����cǎ6�OH��=�����;�i��dLKgʔx��7x��{��ͦ���ꠠ.""҅dd����צ�III���KfF��5�����/�d�޽Xm6RSS����z�d���U�6���kx��o��/��<2o���'����tg�/y.����4h��C�C{�$<x*��?�߆۸���tF;w�d�����`0����j��ҺKK��4҅�n�'� 3#���?����W��QUU�����vS^^���X��=Hjj�w��:s�v;i�i,����ѣ�?�IIIm����EZZ+V�8bd���]?�))):��f����,��7O���=�����H���Ӧr?���HO��O�3�ᇏ�=����������?W�`��������:f�����Ӈ��?k׶�7�E�����<Ì�Ӊ���`0p�m�8眳u�`�KA]DD$B8�����ILH��+�����?=�~������|���Nj��X��csx��̘>�A��p8BӒz�f��˩����S��=**�����5k&/��O>�8��|��C�C{d�s$�`�� >�6ܮ&�6�.i���L�8�]���~jjj��
�V�}�<����9����1j�HRSSy�Y�pa��m2��Z,2��S��"Ȏ��p"/��/-X�ۮs黭��noS9�݁ٔ�Ѻ����_DDD�{999�>��o�b�ٸ�_2fL�n 's�y��O��φذa�o���n��:��/W�ۮs�s�K����Zԛ�y�E�oI-�""�}��u���Rf�y'55�<2��5���r�~�֮�
��Nj��o�����ЮP��������m�fq��]��wW��hQo5ꋡU0o�ݸ4ꋈ�te�sԗC���>l8A�\��������Ķm��z����#F9Y���\v���BZ��κ�:���:tĨ/�CO�����EDD$2�!C��3�P[[�����'Й�]�R���1�z����t&k�~�:h�U�.x<��EDDD �:h�U�������H'3jԨ�-{ʔT�n��u.E��PP��n��������Θ>�;��3ס+��K�y<�M7<9�H��h���yf�|֮�긷H?����!C�2��<�t�:t���s)�u���EDD:aP���A]]_DDDDD"���������������(������(������HG1kD�&����*�jk�x=x<�~X�e2��Z�X-Vbbc���W,������z���POQ���꾳u��~���hjj������=D��&=-�=z蠈���(�w_�`�ݻٿ��� �����E|\<���
�����DuU%�U�����^����o蝔DfF�AIDDDDA�{��|�ع���:�F#}��ЧO*f���p�p8��_f_JJ�QRRL ˶�/+������٘L&,�.������ϰb�
������w����:���i���L!�� ۶�RWW��jeР!�n�2ض-�����ѣ���`0�:d�"�Τ�v�b��ܹ��� ��O<ުܛo�ų�=w�e�u�Ϙ<i o��6�z�}��^/^Lў�#��:t�:������������eKCy�C3ݙ�ٽ����:�V+ÆowH�rF1��a��1�p�����9ݟ{��r�*�6��7X-�V�L��!���7\r�%�y�|����f�ְ��Vu��uضm��_�9]u�8���ٿ���Ƞ�!X���^��jc�!�n���������am)��}�,z��DEE1s�,��):n��Ç�؟�x��i�i�[��뮽��+W����1�=U:_�����܇q8���͚5kU�0�-ꍍ�\4&��s�o��19,|���d�w�1������������O����OyzDG���'���{p�E�����,Y����6QSSÒ%K���׎��EGG���$/7�+���䫯�ٳY�dI���S��r5q�U�x��7��=����y�QJKK����o����ZFu�8Ӣ��?����OqI1��ؘ�328���qӍ7��>��s���+ |�чGt�0��\p��8�=zp�瓖���h�\M���a6�IN��IeYi�F��������8�"]�G}���9n������HLL$&&��Bbb"N�S;0�9��8NJKK���F^�6v����ٳ���ᙧ���������8@u8��y�V�XɴiS��y���_�������O?�o�	�e�P^QAyE�����X�V�����[>?ї�`0xJ�''�y���* ���X,�?-��=��(�1���ܹ���Sg49��C?�|.�����g�؜P�aqq1w��s�+*�绋�5kV�/Z�z�RT�#��_���3�����m�Gu�BA��?`�ȑ��w�%::���Fv��Aa��gͺ�;w�~�p� 0n�X~x.�`���{�E�ޣ���`��Ә8q"S�L	�/���lڼ����\wݵ,X�2�������8p�Q�q��������� �?@��}�6m*�\rI���~vWh��?����@m��on��Occb���jj飠.�e�?.�|߾b��f g�y&i���iEEE��hn!LKM%333�H��_R[[CLL,YY��ر��CbBC������;w�v{�����3�T�|������rJJ
�F�b�e��~�+*���PT���/(����}�v&M� ���>i��L�2��3oU�bPwFEQYUŁu�ڵ����t:1b#F���߿?555�WT4���` ==�'��g�z�m 0���ڕ�SO=͎�;�կ�?�����KbB�qGZy��gx���8k��&�ׯ��̥���]-�-�=�C):�a���=�׍�t-/�2�U�h0�����{ws��f�`4P� yyy���1b��V�lh�gӦ͘�&~?eee444P__��l���QYY���[8��:a�`�.��"���4��_��9�M�NLTT�v|�{�E�=��r��yU���g�:������ܹ��w���HFF:�sS�L	2��sZ�Q�?�����������y�f����hd�܇Y��,]��i7Nc���������&O�L 8�H)eee�n9�f���sɡ������k�����e�t�?��f��}����G��"�HSS��4_H�����g���``��M��SR\L߬,bbbB���~�=�\z���_|I]]-���2���L6m�Dqq1�����2�Bg�y�f�=�H�s
����>c s����X�t/�� ��I\\����ϺiS��p8T��u�0~<Əo5�c�?�{��h=�����e�]Fvv6˖}�����~��Ka�n�-[Ƌ/�@�޽�����������.���/��e|�\曭��z��=�<yr�5�h-��/�/}����ݻ�����÷O��`X�Y"�}������+)))�n.��)��PS[�*�;�P���(��jB������b �������r�ٷ��u��z�Pc��[nfŊ����SQ^N||��\s�drrrTա�u�
��&��Q�����ۛ�5�z����<��_��;��+����:<�&$$�k��99�n6-�Ş\s�͊��ESSS�^L
���;���xc%�Z�^;�b4�Z����ƅ���s���><a��'��Ϊ����w�uw�u���������C�r�9g�����9��b��&�����r��z0d�ҥL�0���ҥ�B��8�V�m��,g��h$ŏ��д��>��s���O.�Zl��\��k�
��ԅ��Y�E����X�ok����>}�`0Z�b�l����DpP߼eK�.��
�N����1��Y}���Ϝu�����K���y뭷Y�z7�0��Lii) �]zi�n/m���̔n��7��ߋ���KZZ���SPXHbbb��_�#&6�ںZ�JKHK�ر��JK�z�bb���F���޽���
>�t9������II���0��;X�r%[s�RYYIcc=��6l�f�ju稜1c�暫�l�g���S^^θ�q �������,-ZD��B�A�߿�_~9ӦN=�������ח�����w�o_1���{�9�sD����ߓ��=�����x:����qs��G�;����;H��2d���Q_� ��у��T�23��DD:��@v;;[<����v5iO4uڍs�E��}�����Juu5QQ=8묑�֯����bcb�<D\D��ŋ��o��罹��]���������̦l��j�m~�8XdŊ��y�O).n�y��yތ�LL&3ee%TTV��TTT���,�Ü��g蠋������zٕ���7n$11�Y3o��+�l�Ng��z�#&��W����ᤷ����ϿX�<�Y�$%%��HDDD$���c歷2�֓��lfF��&~?K�.a̘�m:����*>[���^=1�3�y�=�Pk������zwa080�;��|�'��ۗ3�?����-�7�_�ORrfsxkLLfcНED���8���;^���7�n�d2��=�={
1�L����s�NRR�H�� 6&��Q\����h�n���Kt�hRSS�t�HJJ"##3�'��HW�0F�-�E��PP��of��}��;���"��*��?�WkW��x�z} X,f�V+��Ѥ���ut�����."�n^�����(�w-��A��q�\T�TQWS�����q��²N�Ɉ�b�j�K|\�6-$""Gr���l����(�wIv��>�)�IN���$��@����¦F���%���f���rtU���H���f�d2��r��z�SD�	��CcSc�,KA]DD$A�n�c:�?����˥#�Ź]n��:l�u}	SX�X,��~�~?�MM��l6V�Y���t��ׇ��&�c0B_��EDD"��h��p ��zC���jB��"]��l�d2a�X"#�8Ѐ�jݴADD��Ʉ��$�r�p�ݺɑHu�������/uu���%%���L!�~񈈈|ۡ�\8�N���H���g�����������JA9]DD���""-��;���/+V|�ɨbDD�k�8q�v�����hb��5���-��I�<��������d�E�/�oذ���1�EDDDD��`4��W�ƍy���`�_��q�f�������H��~u������y��4xģ� +V��9g����Ӟ9����5�7��G87|+�7?vH�`n���T�P�c0M��5p۬�9�m����D�6����}�8�g�Qa]DDDD��)�h$����ͮ]{���O2�;�/_��K�c55��Lf���8��ocŊ��4�Iu�1W�ZǅLe�W[�Xm�;������t7�����5�8o�u|���6d�S
���{�s#7N����b��0�-������l""""��by(���6�v�e����؜�(,�w�p�ji����o� s��#G�ɤ�3f�9��HZZ���:�""""�e��7�wo	%%�|��Z�[�_��(��p��:,��%��5���p��'(�ـ`�|���7@DDDD�{����
�-��ўs��.""""ҝ�y[~KP?V@W������(��'��!�-�+�������L66�#��EDDDD����&""""ҝ鶡�%��6"""��� &H�u0u����Q7���<�    IEND�B`�