<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Lägg till ett konto</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="accounts.html" title="Nätkonton">Nätkonton</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Lägg till ett konto</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du lägger till ett konto kommer det bli enklare att länka dina nätkonton med ditt Ubuntu-skrivbord. Din e-post, chattprogram, och andra relaterade program kommer därmed att vara konfigurerade för dig.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ikonen längst till höger i <span class="gui">menyraden</span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Onlinekonton</span>.</p></li>
<li class="steps">
<p class="p">Välj en <span class="gui">kontotyp</span> från fönstrets högra del.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du vill ställa in fler konton kan du upprepa processen när som helst.</p></div></div></div></div>
</li>
<li class="steps"><p class="p">En litet webbgränssnitt kommer öppnas där du kan skriva in uppgifterna för dina nätkonton. Om du till exempel vill lägga till ett Google-konto, skriv in ditt Google-användarnamn, -lösenord, och logga in.</p></li>
<li class="steps"><p class="p">Om du skrev in dina uppgifter korrekt, kommer du tillfrågas om att godkänna villkoren. Välj <span class="gui">Acceptera</span> för att fortsätta. När du har gjort det, behöver Ubuntu tillstånd att komma åt ditt konto. För att ge detta tillstånd, klicka på knappen <span class="gui">Ge åtkomst</span>. När du tillfrågas, skriv in den aktuella användarens lösenord.</p></li>
<li class="steps"><p class="p">Nu kan du välja vilka program du vill länka till ditt onlinekonto. Om du till exempel vill använda ett onlinekonto för chatt, men inte för kalendern, stäng av alternativet <span class="gui">kalender</span>.</p></li>
</ol></div></div></div>
<p class="p">Efter att du har lagt till kontona, kommer alla program du valt automatiskt använda uppgifterna när du loggar in på ditt konto.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Av säkerhetsskäl kommer Ubuntu inte lagra ditt lösenord på din dator. Istället lagras en slags bricka som kommer från onlinetjänsten. Om du vill återkalla länken mellan ditt skrivbord och onlinetjänsten, <span class="link"><a href="accounts-remove.html" title="Ta bort ett konto">ta bort</a></span> den.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="accounts.html" title="Nätkonton">Nätkonton</a><span class="desc"> — <span class="link"><a href="accounts-add.html" title="Lägg till ett konto">Lägg till kontakter, </a></span> <span class="link"><a href="accounts-remove.html" title="Ta bort ett konto">Ta bort konton, </a></span> <span class="link"><a href="accounts-disable-service.html" title="Avaktivera kontotjänster">Avaktivera tjänster</a></span></span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
