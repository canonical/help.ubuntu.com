<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vad är nytt i Ubuntu 14.04?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Vad är nytt i Ubuntu 14.04?</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Med Ubuntu 14.04 LTS fortsätter utvecklingen av <span class="em">Unity</span>-gränssnittet. Nedan finner du några av de viktigaste förändringarna sedan Ubuntu 12.04 LTS.</p></div>
<div id="new-features" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Nya och förbättrade funktioner</span></h2></div>
<div class="region"><div class="contents"><div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Menyerna till det program som är i fokus är som standard tillgängliga på Ubuntus integrerade <span class="link"><a href="unity-menubar-intro.html#app-menus" title="Programmenyer">menylist</a></span>. Du kan dock byta till den konventionella stilen, om du vill, och visa programmenyerna på namnlisten i fönstret för respektive program i stället (den senare möjligheten är ny sedan Ubuntu 13.10).</p></li>
<li class="list"><p class="p">Det har tillkommit stöd för att ändra Unitys skärmupplösning separat för varje ansluten monitor, vilket gör det lättare att använda skärmar med hög upplösning. Liknande stöd finns även i LibreOffice och Chromium.</p></li>
<li class="list"><p class="p">Förbättrat utseende såsom rundade fönsterdekorationer, ett nytt gränssnitt för att låsa upp skärmen, och andra stiljusteringar.</p></li>
<li class="list"><p class="p">Det <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">integrerade <span class="gui">Textinmatning</span>s-gränssnittet</a></span> och den tillhörande <span class="link"><a href="unity-menubar-intro.html#status-menus" title="Statusmenyer">indikatorn</a></span> för inmatningskällor är utformade för att ställa in både tangentbordslayout och IBus-inmatningsmetoder.</p></li>
<li class="list">
<p class="p"><span class="gui">Dash</span> har genomgått ett antal förbättringar:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p"><span class="gui">Dash</span> kan nu söka bland dussintals källor på Internet samtidigt. Funktionen att söka på Internet <span class="link"><a href="unity-shopping.html" title="Varför finns det shoppinglänkar i Dash?">kan inaktiveras</a></span>.</p></li>
<li class="list"><p class="p">Sökresultaten från <span class="gui">Dash</span> kan filtreras per kategori och källa..</p></li>
<li class="list"><p class="p">Genom att högerklicka på ett sökresultat i <span class="gui">Dash</span> visas en ruta med förhandsinformation.</p></li>
<li class="list"><p class="p">Använd <span class="link"><a href="unity-dash-photos.html" title="Fotolinsen">fotolinsen</a></span> för att se foton på datorn eller på dina konton i sociala medier.</p></li>
<li class="list"><p class="p">Anpassa <span class="gui">Dash</span> genom att lägga till och ta bort linser.</p></li>
<li class="list"><p class="p">Läs meddelanden från dina konton på sociala medier genom den nya funktionen <span class="link"><a href="unity-dash-friends.html" title="Vänner">Vänner</a></span>.</p></li>
</ul></div></div></div>
</li>
<li class="list"><p class="p">Ange dina inloggingsuppgifter i <span class="link"><a href="accounts.html" title="Nätkonton">Nätkonton</a></span> för att enkelt sätta upp samordning för till exempel Dash och Empathy.</p></li>
<li class="list"><p class="p">Håll reda på kontaktuppgifter till dina vänner och kollegor genom <span class="link"><a href="contacts.html" title="Kontakter">Kontakter</a></span>, din personliga adressbok.</p></li>
</ul></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links ">
<a href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord, program &amp; fönster</a><span class="desc"> — <span class="link"><a href="unity-introduction.html" title="Välkommen till Ubuntu">Introduktion</a></span>, <span class="link"><a href="shell-keyboard-shortcuts.html" title="Användbara kortkommandon">kortkommandon</a></span>, <span class="link"><a href="shell-windows.html" title="Fönster och arbetsytor">fönster</a></span>…</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
