<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använd andra högtalar eller hörlurar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="media.html#sound" title="Grundinställningar ljud">Ljud</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Använd andra högtalar eller hörlurar</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan använda externa högtalare eller hörlurar med din dator. Högtalare kopplas vanligtvis via en cirkulär teleplugg eller via USB.</p>
<p class="p">Om dina högtalare eller hörlurar har en teleplugg, koppla in den i en lämplig kontakt på din dator. De flesta datorer har två kontakter: en för mikrofoner och en för högtalare. Leta efter en bild på hörlurar intill kontakten. Högtalare eller hörlurar som kopplats in i en telepluggskontakt kommer vanligtvis att användas som standard. Om inte, se instruktionerna nedan för att välja standardenheten.</p>
<p class="p">Vissa datorer har stöd för flerkanalsutmatning för surround-ljud. Detta kräver i regel flera TRS-jack, som oftast är färgkodade. Om du inte är säker på vilka kontakter sladdarna ska sitta i kan du testa ljudutmatningen i ljudinställningarna. Klicka på <span class="gui">ljudmenyn</span> på <span class="gui">menyraden</span> och klicka sedan på <span class="gui">Ljudinställningar</span>. Välj dina högtalare i listan över enheter, och klicka sedan på <span class="gui">Testa ljud</span>. I fönstret som dyker upp, klicka på knappen för varje högtalare. Varje knapp bör läsa upp sin position endast i den kanal som motsvarar den högtalaren.</p>
<p class="p">Om du har USB-högtalare eller hörlurar eller analoga hörlurar kopplade i ett USB-ljudkort kan du koppla in dem i vilken USB-kontakt som helst. USB-högtalare fungerar som separata ljudenheter och du kan behöver ange vilka högtalar som ska användas som standard.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Välj en standard ljudinmatningsenhet</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="gui">ljudmenyn</span> på <span class="gui">menyraden</span> och välj <span class="gui">Ljudinställningar</span>.</p></li>
<li class="steps"><p class="p">På fliken <span class="gui">Utmatning</span>, välj enheten i listan.</p></li>
</ol></div>
</div></div>
<p class="p">Om du inte ser din enhet på fliken <span class="gui">Utmatning</span>, kontrollera fliken <span class="gui">Hårdvara</span>. Välj din enhet och testa olika profiler.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="media.html#sound" title="Grundinställningar ljud">Grundinställningar ljud</a><span class="desc"> — <span class="link"><a href="sound-volume.html" title="Ändra ljudvolymen">Volym</a></span>, <span class="link"><a href="sound-usespeakers.html" title="Använd andra högtalar eller hörlurar">högtalare och hörlurar</a></span>, <span class="link"><a href="sound-usemic.html" title="Använd en annan mikrofon">mikrofoner</a></span>...</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="sound-usemic.html" title="Använd en annan mikrofon">Använd en annan mikrofon</a><span class="desc"> — Använd en analog eller USB-mikrofon och välj standardingångsenhet.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
