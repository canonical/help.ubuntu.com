<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Hitta program, filer, musik och annat med Dash</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Hitta program, filer, musik och annat med Dash</span></h1></div>
<div class="region">
<div class="contents">
<div class="media media-image floatend"><div class="inner"><img src="figures/unity-dash-sample.png" class="media media-block" alt="Unity Search"></div></div>
<p class="p">The <span class="gui">Dash</span> allows you to search for applications, files, music, and videos,
    and shows you items that you have used recently. If you have ever worked on
    a spreadsheet or edited an
    image and forgot where you saved it, you will surely find this feature of the Dash to be useful.
  </p>
<p class="p">To start using the <span class="gui">Dash</span>, click the top icon in the <span class="link"><a href="unity-launcher-intro.html" title="Använda programstartaren">Launcher</a></span>.
    This icon has the Ubuntu logo on it.
    For faster access, you can just press the <span class="key"><a href="windows-key.html" title='Vad är "Superknappen"?'><kbd>Super</kbd></a></span> key.</p>
<p class="p">To hide the <span class="gui">Dash</span>, click the top icon again or press <span class="key"><kbd>Super</kbd></span> or <span class="key"><kbd>Esc</kbd></span>.</p>
</div>
<div id="dash-home" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Search everything from the Dash home</span></h2></div>
<div class="region">
<div class="contents">
<p class="p">The first thing you'll see when opening the Dash is the Dash Home. Without typing
    or clicking anything, the Dash Home will show you apps and files you've used recently.</p>
<p class="p">Only one row of results will show for each type. If there are more results, you can
    click <span class="gui">See more results</span> to view them.</p>
<p class="p">To search, just start typing and related search results will automatically appear
    from the different installed lenses.</p>
<p class="p">Click on a result to open it, or you can press <span class="key"><kbd>Enter</kbd></span> to open the first
    item in the list.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="shell-apps-favorites.html" title="Change which applications show in the Launcher">Change which applications show in the Launcher</a><span class="desc"> — Add, move, or remove frequently-used program icons on the 
    Launcher.</span>
</li>
<li class="links ">
<a href="unity-shopping.html" title="Varför finns det shoppinglänkar i Dash?">Varför finns det shoppinglänkar i Dash?</a><span class="desc"> — Online results make the Dash more useful and help fund Ubuntu 
    development.</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="dash-lenses" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Lenses</span></h2></div>
<div class="region">
<div class="contents">
<p class="p">Lenses allow you to focus the Dash results and exclude results from other lenses.</p>
<p class="p">You can see the available lenses in the <span class="gui">lens bar</span>, the darker strip at
    the bottom of the Dash.</p>
<p class="p">To switch to a different lens, click the appropriate icon or press
    <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span>.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="unity-dash-apps.html" title="Applications lens">Applications lens</a><span class="desc"> — Run, install, or uninstall apps.</span>
</li>
<li class="links ">
<a href="unity-dash-files.html" title="Files lens">Files lens</a><span class="desc"> — Find files, folders, and downloads.</span>
</li>
<li class="links ">
<a href="unity-dash-photos.html" title="Fotolinsen">Fotolinsen</a><span class="desc"> — View photos from your computer or your online social media 
    accounts.</span>
</li>
<li class="links ">
<a href="unity-dash-music.html" title="Music lens">Music lens</a><span class="desc"> — Find and play music from your computer or the internet.</span>
</li>
<li class="links ">
<a href="unity-dash-video.html" title="Video lens">Video lens</a><span class="desc"> — Find and play videos from your computer or the internet.</span>
</li>
<li class="links ">
<a href="unity-dash-friends.html" title="Vänner">Vänner</a><span class="desc"> — Browse messages from your online social media accounts.</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="dash-filters" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Filters</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Filters allow you to narrow down your search even further.</p>
<p class="p">Click <span class="gui">Filter results</span> to choose filters. You may need to click a
    filter heading such as <span class="gui">Sources</span> to see the available choices.</p>
</div></div>
</div></div>
<div id="dash-previews" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Previews</span></h2></div>
<div class="region"><div class="contents">
<p class="p">If you right click on a search result, a <span class="gui">preview</span> will open with more
    information about the result.</p>
<p class="p">To close the preview, click any empty space or press <span class="key"><kbd>Esc</kbd></span>.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
