<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Växla uppgifter</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 21.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="getting-started.html.sv" title="Komma igång">Kom igång med GNOME</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<nav class="prevnext pagewide"><div class="inner">
<a href="gs-launch-applications.html.sv" title="Starta program">Föregående</a><a href="gs-use-windows-workspaces.html.sv" title="Använda fönster och arbetsytor">Nästa</a>
</div></nav><div class="hgroup pagewide"><h1 class="title"><span class="title">Växla uppgifter</span></h1></div>
<div class="region">
<div class="contents pagewide"><div class="links-tile">
<a href="figures/gnome-task-switching.webm" class="ui-overlay"><span class="links-tile-img"><img src="gs-thumb-task-switching.svg" width="812"></span></a><div class="ui-overlay"><div class="inner">
<a href="#" class="ui-overlay-close" title="Stäng">⨯</a><div class="contents"><div class="media media-video"><div class="inner">
<video src="figures/gnome-task-switching.webm" preload="auto" class="media media-block" height="394" width="700"></video><div class="media-controls media-controls-video media-controls-ttml">
<button class="media-play" data-play-label="Spela upp" data-pause-label="Paus" value="Spela upp"><svg width="20" height="20" class="media-play"><polygon points="5,4 5,16 15,10" class="yelp-svg-fill"></polygon></svg><svg width="20" height="20" class="media-pause"><rect x="4" y="4" width="4" height="12" class="yelp-svg-fill"></rect><rect x="12" y="4" width="4" height="12" class="yelp-svg-fill"></rect></svg></button><input type="range" class="media-range" value="0"><span class="media-time"><span class="media-current">0:00</span><span class="media-duration">-:--</span></span>
</div>
<div class="media-ttml">
<div class="media-ttml-node media-ttml-div" data-ttml-begin="1" data-ttml-end="5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="1" data-ttml-end="5">Växlar uppgifter</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="5" data-ttml-end="8"><div class="media-ttml-node media-ttml-p" data-ttml-begin="5" data-ttml-end="8">Flytta din musmarkör till <span class="gui">Aktivitetshörnet</span> längst upp till vänster på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="9" data-ttml-end="12"><div class="media-ttml-node media-ttml-p" data-ttml-begin="9" data-ttml-end="12">Klicka på ett fönster för att byta till den uppgiften.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="12" data-ttml-end="14"><div class="media-ttml-node media-ttml-p" data-ttml-begin="12" data-ttml-end="14">För att maximera ett fönster längs skärmens vänstra sida, fånga fönstrets namnlist och dra det åt vänster.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="14" data-ttml-end="16"><div class="media-ttml-node media-ttml-p" data-ttml-begin="14" data-ttml-end="16">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="16" data-ttml-end="0"><div class="media-ttml-node media-ttml-p" data-ttml-begin="16" data-ttml-end="0">För att maximera ett fönster längs den högra sidan, fånga fönstrets namnlist och dra det åt höger.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="18" data-ttml-end="20"><div class="media-ttml-node media-ttml-p" data-ttml-begin="18" data-ttml-end="20">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="23" data-ttml-end="27"><div class="media-ttml-node media-ttml-p" data-ttml-begin="23" data-ttml-end="27">Tryck <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>+<span class="key"><kbd> Tabb</kbd></span></span> för att visa <span class="gui">fönsterväxlaren</span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="27" data-ttml-end="29"><div class="media-ttml-node media-ttml-p" data-ttml-begin="27" data-ttml-end="29">Släpp <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> för att välja nästa markerade fönster.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="29" data-ttml-end="32"><div class="media-ttml-node media-ttml-p" data-ttml-begin="29" data-ttml-end="32">För att bläddra igenom listan av öppna fönster, släpp inte <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> utan håll den nertryckt och tryck på <span class="key"><kbd>Tabb</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="35" data-ttml-end="37"><div class="media-ttml-node media-ttml-p" data-ttml-begin="35" data-ttml-end="37">Tryck på <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super </kbd></a></span> för att visa <span class="gui">Aktivitetsöversikt</span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="37" data-ttml-end="40"><div class="media-ttml-node media-ttml-p" data-ttml-begin="37" data-ttml-end="40">Börja skriv in namnet på det program du vill växla till.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="40" data-ttml-end="43"><div class="media-ttml-node media-ttml-p" data-ttml-begin="40" data-ttml-end="43">När programmet visas som det första resultatet, tryck på <span class="key"><kbd>Retur</kbd></span> för att växla till det.</div></div>
</div>
</div></div></div>
</div></div>
</div></div>
<section id="switch-tasks-overview"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Växla uppgifter</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Flytta din musmarkör till <span class="gui">Aktiviteter</span>-hörnet längst upp till vänster på skärmen för att via <span class="gui">Aktivitetsöversikt</span> där du kan se alla de körande uppgifterna visas som små fönster.</p></li>
<li class="steps"><p class="p">Klicka på ett fönster för att byta till den uppgiften.</p></li>
</ol></div></div></div></div></div>
</div></section><section id="switching-tasks-tiling"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Lägg fönster sida-vid-sida</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">För att maximera ett fönster längs en sida av skärmen, fånga fönstrets namnlist och dra det till vänster eller höger sida av skärmen.</p></li>
<li class="steps"><p class="p">När hälften av skärmen är markerad, släpp fönstret för att maximera det längs den valda sidan av skärmen.</p></li>
<li class="steps"><p class="p">För att maximera två fönster sida-vid-sida, fånga namnlisten på det andra fönstret och dra det till den andra sidan av skärmen.</p></li>
<li class="steps"><p class="p">När hälften av skärmen är markerad, släpp fönstret för att maximera det längs den andra sidan av skärmen.</p></li>
</ol></div></div></div></div></div>
</div></section><section id="switch-tasks-windows"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Växla mellan fönster</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Tryck på <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super </kbd></a></span>+<span class="key"><kbd>Tabb</kbd></span></span> för att visa <span class="gui">fönsterväxlaren</span>, som listar alla öppna fönster.</p></li>
<li class="steps"><p class="p">Släpp <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> för att välja nästa markerade fönster i <span class="gui">fönsterväxlaren</span>.</p></li>
<li class="steps"><p class="p">För att bläddra igenom listan av öppna fönster, släpp inte <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> utan håll den nertryckt och tryck på <span class="key"><kbd>Tabb</kbd></span>.</p></li>
</ol></div></div></div></div></div>
</div></section><section id="switch-tasks-search"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Använd sökning för att växla mellan program</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Tryck på <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> för att visa <span class="gui">Aktivitetsöversikt</span>.</p></li>
<li class="steps"><p class="p">Bara börja skriv namnet på det program du vill växla till. Program som matchar det du har skrivit kommer att visas medan du skriver.</p></li>
<li class="steps"><p class="p">När programmet som du vill växla till visas som det första resultatet, tryck på <span class="key"><kbd>Retur</kbd></span> för att växla till det.</p></li>
</ol></div></div></div></div></div>
</div></section><nav class="prevnext pagewide"><div class="inner">
<a href="gs-launch-applications.html.sv" title="Starta program">Föregående</a><a href="gs-use-windows-workspaces.html.sv" title="Använda fönster och arbetsytor">Nästa</a>
</div></nav><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="getting-started.html.sv" title="Komma igång">Kom igång med GNOME</a><span class="desc"> — Är GNOME nytt för dig? Lär dig hur du använder det.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-windows-switching.html.sv" title="Växla mellan fönster">Växla mellan fönster</a><span class="desc"> — Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span>.</span>
</li></ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
