<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>dpkg</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = "index.html.en";
        } else {
                window.location = href.replace(/\.html.*/, ".html.en");
        }
         return false;
      }
      function browserPreferredLanguage() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = href;
        } else {
                window.location = href.replace(/\.html.*/, ".html");
        }
        return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../18.04" class="trail">Ubuntu 18.04</a> » <a class="trail" href="index.html.sv" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="package-management.html.sv" title="Pakethantering">Pakethantering</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="package-management-introduction.html.sv" title="Inledning">Föregående</a><a class="nextlinks-next" href="apt.html.sv" title="Apt">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">dpkg</h1></div>
<div class="region"><div class="contents">
<p class="para">
    <span class="app application">dpkg</span> is a package manager for <span class="em emphasis">Debian</span>-based systems.  It can install, remove, and build packages, but
    unlike other package management systems, it cannot automatically download and install packages or their dependencies.  This section covers using
    <span class="app application">dpkg</span> to manage locally installed packages:
    </p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">

        <p class="para">
        To list all packages installed on the system, from a terminal prompt type:
        </p>

<div class="screen"><pre class="contents "><span class="cmd command">dpkg -l</span>
</pre></div>

      </li>
<li class="list itemizedlist">

        <p class="para">Beroende på mängden paket i ditt system, så kan det generera en stor mängd utdata.  Rikta utdatan genom <span class="app application">grep</span> för att se om ett specifikt paket är installerat:</p>

<div class="screen"><pre class="contents "><span class="cmd command">dpkg -l | grep apache2</span>
</pre></div>

        <p class="para">Ersätt <span class="em emphasis">apache2</span> med något paketnamn, del av paketnamn eller annat reguljärt uttryck.</p>

      </li>
<li class="list itemizedlist">

        <p class="para">För att lista filer som installerats av ett paket, i det här fallet paketet <span class="app application">ufw</span>, skriv:</p>

<div class="screen"><pre class="contents "><span class="cmd command">dpkg -L ufw</span>
</pre></div>

      </li>
<li class="list itemizedlist">

        <p class="para">Om du är osäker på vilket paket som installerat en fil, då kan kanske <span class="app application">dpkg -S</span> ge dig en förklaring. Till exempel:</p>

<div class="screen"><pre class="contents "><span class="cmd command">dpkg -S /etc/host.conf</span>
<span class="output computeroutput">base-files: /etc/host.conf</span>
</pre></div>

        <p class="para">Resultatet visar att <span class="file filename">/etc/host.conf</span> tillhör paketet <span class="app application">base-files</span>.</p>

        <div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
          <p class="para">
          Many files are automatically generated during the package install process, and even though they are on the filesystem, 
          <span class="cmd command">dpkg -S</span> may not know which package they belong to.
          </p>
        </div></div></div></div>

      </li>
<li class="list itemizedlist">

        <p class="para">Du kan installera en lokal <span class="em emphasis">.deb</span>-fil genom att skriva:</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo dpkg -i zip_3.0-4_i386.deb</span>
</pre></div>
    
        <p class="para">
        Change <span class="file filename">zip_3.0-4_i386.deb</span> to the actual file name of the local .deb file you wish to install.
        </p>

      </li>
<li class="list itemizedlist">

        <p class="para">Avinstallera ett paket verkställs genom:</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo dpkg -r zip</span>
</pre></div>

        <div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents">
          <p class="para">
          Uninstalling packages using <span class="app application">dpkg</span>, in most cases, is <span class="em emphasis">NOT</span> recommended.
          It is better to use a package manager that handles dependencies to ensure that the system is in a consistent state.  For
          example using <span class="cmd command">dpkg -r zip</span> will remove the <span class="app application">zip</span> package, but any packages that
          depend on it will still be installed and may no longer function correctly.
          </p>
        </div></div></div></div>

      </li>
</ul></div>
<p class="para">För fler alternativ till <span class="app application">dpkg</span> se manualsidan: <span class="cmd command">man dpkg</span>.</p>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="package-management-introduction.html.sv" title="Inledning">Föregående</a><a class="nextlinks-next" href="apt.html.sv" title="Apt">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address
          so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>
          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p>
</div>
</div>
</body>
</html>
