<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Dela ut och överför filer</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="sharing.html" title="Sharing">Sharing</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Dela ut och överför filer</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan dela filer med dina kontakter, eller överföra dem till externa enheter eller <span class="link"><a href="nautilus-connect.html" title="Bläddra bland filer på en server eller nätverksdelning">nätverksdelningar</a></span> direkt från filhanteraren.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna <span class="link"><a href="files-browse.html" title="Bläddra bland filer och mappar">filhanteraren</a></span>.</p></li>
<li class="steps"><p class="p">Hitta filen du vill överföra.</p></li>
<li class="steps"><p class="p">Högerklicka på filen och välj <span class="gui">Skicka till</span>.</p></li>
<li class="steps"><p class="p">Fönstret <span class="gui">Skicka till</span> kommer visas. Välj vart du vill skicka filen och klicka på <span class="gui">Skicka</span>. Se listan över destinationer nedanför för mer information.</p></li>
</ol></div></div></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan skicka flera filer vid samma tillfälle. Markera flera filer genom att hålla ner <span class="key"><kbd>Ctrl</kbd></span>, och högerklicka sedan på en av de markerade filerna. Du kan automatiskt komprimera filerna till ett zip- eller tar-arkiv.</p></div></div></div></div>
<div class="list"><div class="inner">
<div class="title title-list"><h2><span class="title">Mål</span></h2></div>
<div class="region"><ul class="list">
<li class="list"><p class="p">För att e-posta filen, välj <span class="gui">E-post</span> och skriv in mottagarens e-postadress.</p></li>
<li class="list"><p class="p">För att skicka filen till en snabbmeddelandeklient, välj <span class="gui">Snabbmeddelande</span> och välj sedan en kontakt från den utfällbara listan. Ditt snabbmeddelandeprogram kan behöva ha startats för att det ska fungera.</p></li>
<li class="list"><p class="p">För att bränna filerna till en cd- eller dvd-skiva, välj <span class="gui">cd-/dvd-skaparen</span>. Se <span class="link"><a href="files-disc-write.html" title="Skriv filer till en cd- eller dvd-skiva">Skriv filer till en cd- eller dvd-skiva</a></span> för mer information.</p></li>
<li class="list"><p class="p">För att föra över filen till en Bluetooth-enhet, välj <span class="gui">Bluetooth (OBEX Push)</span> och välj enheten du vill skicka filen till. Du kommer bara se enheter du redan har parat med. Se <span class="link"><a href="bluetooth.html" title="Bluetooth">Bluetooth</a></span> för mer information.</p></li>
<li class="list"><p class="p">För att kopiera en fil till en extern enhet, som ett USB-minne, eller ladda upp den till en server du är ansluten till, välj <span class="gui">Flyttbara diskar och delningar</span>, och välj sedan enheten eller servern du vill kopiera filen till.</p></li>
</ul></div>
</div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li>
<li class="links ">
<a href="sharing.html" title="Sharing">Sharing</a><span class="desc"> — 
      <span class="link"><a href="sharing-desktop.html" title="Share your desktop">Desktop sharing</a></span>,
      <span class="link"><a href="files-share.html" title="Dela ut och överför filer">Share files</a></span>…
    </span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="nautilus-connect.html" title="Bläddra bland filer på en server eller nätverksdelning">Bläddra bland filer på en server eller nätverksdelning</a><span class="desc"> — Visa och redigera filer på en annan dator över FTP, SSH, Windows-delningar, eller WebDAV.</span>
</li>
<li class="links ">
<a href="bluetooth-send-file.html" title="Skicka en fil till en Bluetooth-enhet">Skicka en fil till en Bluetooth-enhet</a><span class="desc"> — Dela filer till Bluetooth-enheter som din telefon.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
