<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Inställningar för användare och system</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Inställningar för användare och system</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-grid ">
<div class="links-grid-link"><a href="user-accounts.html" title="Användarkonton">Användarkonton</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="user-add.html" title="Lägg till ett nytt användarkonto">Lägg till användare</a></span>, <span class="link"><a href="user-changepassword.html" title="Välj ditt lösenord">ändra lösenord</a></span>, <span class="link"><a href="user-admin-change.html" title="Ändra vem som har administratörsbehörighet">administratörer</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="clock.html" title="Datum och tid">Datum och tid</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="clock-set.html" title="Ändra datum och tid">Sätt datum och tid</a></span>, <span class="link"><a href="clock-world.html" title="Lägg till en världsklocka">världsklockor</a></span>, <span class="link"><a href="clock-timezone.html" title="Ändra din tidszon">tidszon</a></span>, <span class="link"><a href="clock-calendar.html" title="Kalendermöten">kalender och möten</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="prefs-sharing.html" title="Dela-inställningar">Dela-inställningar</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="sharing-bluetooth.html" title="Styr delning över Bluetooth">Bluetooth-delning</a></span>, <span class="link"><a href="sharing-personal.html" title="Dela ut dina personliga filer">Delning av personliga filer</a></span>, <span class="link"><a href="sharing-desktop.html" title="Dela ditt skrivbord">Skärmdelning</a></span>, <span class="link"><a href="sharing-media.html" title="Dela din musik, foton och videor">Mediadelning</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="color.html" title="Färghantering">Färghantering</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="color-whyimportant.html" title="Varför är färghantering viktigt?">Varför är detta viktigt</a></span>, <span class="link"><a href="color.html#profiles" title="Färgprofiler">Färgprofiler</a></span>, <span class="link"><a href="color.html#calibration" title="Kalibrering">Hur du kalibrerar en enhet</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="media.html#sound" title="Grundläggande ljud">Ljud</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="sound-volume.html" title="Ändra ljudvolymen">Volym</a></span>, <span class="link"><a href="sound-usespeakers.html" title="Använd andra högtalar eller hörlurar">högtalare och hörlurar</a></span>, <span class="link"><a href="sound-usemic.html" title="Använd en annan mikrofon">mikrofoner</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="mouse.html" title="Mus">Mus</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="mouse-lefthanded.html" title="Använd din mus med vänster hand">Vänsterhänt</a></span>, <span class="link"><a href="mouse-sensitivity.html" title="Justera hastigheten för musen och styrplattan">hastighet och känslighet</a></span>, <span class="link"><a href="mouse-touchpad-click.html" title="Klicka, dra eller rulla med styrplattan">klickning och rullning med styrplatta</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="accounts.html" title="Nätkonton">Nätkonton</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="accounts-add.html" title="Lägg till ett konto">Lägg till ett nätkonto</a></span>, <span class="link"><a href="accounts-remove.html" title="Ta bort ett konto">Ta bort ett konto</a></span>, <span class="link"><a href="accounts-which-application.html" title="Nättjänster och program">Lär dig om tjänster</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="prefs-language.html" title="Region &amp; språk">Region &amp; språk</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="session-language.html" title="Ändra vilket språk du använder">Ändra språk</a></span>, <span class="link"><a href="session-formats.html" title="Ändra datum och mätvärden">region och format</a></span>, <span class="link"><a href="keyboard-layouts.html" title="Use alternative keyboard layouts">tangentbordslayouter</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="privacy.html" title="Sekretessinställningar">Sekretessinställningar</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="privacy-screen-lock.html" title="Lås automatiskt din skärm">Skärmlås</a></span>, <span class="link"><a href="privacy-history-recent-off.html" title="Stäng av eller begränsa filhistorik">Användningshistorik</a></span>, <span class="link"><a href="privacy-purge.html" title="Töm papperskorgen &amp; ta bort tillfälliga filer">Ta bort skräp &amp; temporära filer</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="power.html" title="Ström och batteri">Ström och batteri</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="power-status.html" title="Kontrollera batteristatus">Batteristatus</a></span>, <span class="link"><a href="power-suspend.html" title="Vad händer när jag försätter min dator i vänteläge?">försätta i vänteläge</a></span>, <span class="link"><a href="power-whydim.html" title="Varför tonas min skärm ner efter ett tag?">skärmtoning</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="keyboard-layouts.html" title="Use alternative keyboard layouts">Tangentbordslayouter</a></span>, <span class="link"><a href="keyboard-cursor-blink.html" title="Få tangentbordsmarkören att blinka">markörblinkning</a></span>, <span class="link"><a href="a11y.html#mobility" title="Rörelsehinder">tangentbordshjälpmedel</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="startup-applications.html" title="Uppstartsprogram">Uppstartsprogram</a></div>
<div class="desc"><span class="desc">Välj vilka program som skall startas när du loggar in.</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="prefs-display.html" title="Visning och skärm">Visning och skärm</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="look-background.html" title="Ändra skrivbords- och låsskärmsbakgrunderna">Bakgrund</a></span>, <span class="link"><a href="look-resolution.html" title="Ändra upplösning eller rotation på skärmen">storlek och rotering</a></span>, ljusstyrka…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="wacom.html" title="Wacom ritplatta">Wacom ritplatta</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="wacom-multi-monitor.html" title="Välj en skärm">Mappa en skärm</a></span>, <span class="link"><a href="wacom-stylus.html" title="Konfigurera pennan">konfigurera pennan</a></span>, <span class="link"><a href="wacom-left-handed.html" title="Använd plattan med vänster hand">använd plattan med vänster hand</a></span>…</span></div>
</div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
