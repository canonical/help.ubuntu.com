<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Utskrifter</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Utskrifter</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="printing-inklevel.html.sv" title="Hur kan jag kontrollera min skrivares bläck- eller tonernivå?"><span class="title">Hur kan jag kontrollera min skrivares bläck- eller tonernivå?</span><span class="linkdiv-dash"> — </span><span class="desc">Kontrollera mängden bläck eller toner som finns kvar i skrivarpatroner.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="printing-to-file.html.sv" title="Skriv ut till fil"><span class="title">Skriv ut till fil</span><span class="linkdiv-dash"> — </span><span class="desc">Spara ett dokument som en PDF-, Postscript- eller SVG-fil istället för att skicka den till en skrivare.</span></a></div>
</div></div></div></div>
<div id="setup" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ställ in en skrivare</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="printing-setup.html.sv" title="Ställ in en lokal skrivare"><span class="title">Ställ in en lokal skrivare</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in en skrivare som är ansluten till din dator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="printing-setup-default-printer.html.sv" title="Ställ in standardskrivaren"><span class="title">Ställ in standardskrivaren</span><span class="linkdiv-dash"> — </span><span class="desc">Välj skrivaren som du använder oftast.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="printing-name-location.html.sv" title="Ändra namnet eller platsen för en skrivare"><span class="title">Ändra namnet eller platsen för en skrivare</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra namnet eller platsen för en skrivare i skrivarinställningarna.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="paper" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Olika pappersstorlekar och layouter</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="printing-select.html.sv" title="Skriv endast ut vissa sidor"><span class="title">Skriv endast ut vissa sidor</span><span class="linkdiv-dash"> — </span><span class="desc">Skriv bara ut specifika sidor, eller ett intervall av sidor.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="printing-2sided.html.sv" title="Skriv ut dubbelsidigt och flersidslayouter"><span class="title">Skriv ut dubbelsidigt och flersidslayouter</span><span class="linkdiv-dash"> — </span><span class="desc">Skriv ut på båda sidorna av pappret eller flera sidor per ark.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="printing-booklet.html.sv" title="Skriv ut ett häfte"><span class="title">Skriv ut ett häfte</span><span class="linkdiv-dash"> — </span><span class="desc">Hur du skriver ut ett vikt, flersidigt häfte med A4 eller papper i Letter-storlek.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="printing-order.html.sv" title="Skriv ut sidor i en annan ordning"><span class="title">Skriv ut sidor i en annan ordning</span><span class="linkdiv-dash"> — </span><span class="desc">Sortera och omvänd utskriftsordningen.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="printing-envelopes.html.sv" title="Skriva ut kuvert"><span class="title">Skriva ut kuvert</span><span class="linkdiv-dash"> — </span><span class="desc">Säkerställ att du har kuvertet med rätt sida upp och har valt den korrekta pappersstorleken.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="printing-differentsize.html.sv" title="Ändra pappers storlek vid utskrift"><span class="title">Ändra pappers storlek vid utskrift</span><span class="linkdiv-dash"> — </span><span class="desc">Skriv ut ett dokument på en annan pappersstorlek eller orientering.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="problems" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Skrivarproblem</span></h2></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="printing-cancel-job.html.sv" title="Avbryt, pausa eller släpp ett utskriftsjobb"><span class="title">Avbryt, pausa eller släpp ett utskriftsjobb</span><span class="linkdiv-dash"> — </span><span class="desc">Hur du avbryter ett väntande jobb och tar bort det från kön.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="printing-paperjam.html.sv" title="Hur du reder ut papperstrassel"><span class="title">Hur du reder ut papperstrassel</span><span class="linkdiv-dash"> — </span><span class="desc">Hur du reder ut papperstrassel beror på tillverkare och modell av skrivaren som du har.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="printing-streaks.html.sv" title="Varför finns det streck, linjer eller fel färger på mina utskrifter?"><span class="title">Varför finns det streck, linjer eller fel färger på mina utskrifter?</span><span class="linkdiv-dash"> — </span><span class="desc">Om utskrifter är streckade, tonande eller saknar färger, kontrollera dina bläcknivåer eller rensa skrivarhuvudet.</span></a></div></div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h3><span class="title">Mer information</span></h3></div>
<div class="region"><ul><li class="links "><a href="hardware.html.sv#problems" title="Vanliga problem">Hårdvaruproblem</a></li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="hardware.html.sv" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a><span class="desc"> — <span class="link"><a href="hardware.html.sv#problems" title="Vanliga problem">Hårdvaruproblem</a></span>, <span class="link"><a href="printing.html.sv" title="Utskrifter">skrivare</a></span>, <span class="link"><a href="power.html.sv" title="Ström och batteri">ströminställningar</a></span>, <span class="link"><a href="color.html.sv" title="Färghantering">färghantering</a></span>, <span class="link"><a href="bluetooth.html.sv" title="Bluetooth">Bluetooth</a></span>, <span class="link"><a href="disk.html.sv" title="Diskar och lagring">diskar</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
