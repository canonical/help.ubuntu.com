<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Filesystem</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="cgroups.html" title="Control Groups">Control Groups</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups-overview.html" title="Översikt">Föregående</a><a class="nextlinks-next" href="cgroups-delegation.html" title="Delegation">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Filesystem</h1></div>
<div class="region"><div class="contents">
<p class="para">
A hierarchy is created by mounting an instance of the cgroup filesystem
with each of the desired subsystems listed as a mount option.  For instance,
  </p>
<div class="screen"><pre class="contents "><span class="cmd command">
mount -t cgroup -o devices,memory,freezer cgroup /cgroup1
</span></pre></div>
<p class="para">
would instantiate a hierarchy with the devices and memory cgroups comounted.
A child cgroup "child1" can be created using 'mkdir'
  </p>
<div class="screen"><pre class="contents "><span class="cmd command">
mkdir /cgroup1/child1
</span></pre></div>
<p class="para">
and tasks can be moved into the new child cgroup by writing their process
IDs into the 'tasks' or 'cgroup.procs' file:
  </p>
<div class="screen"><pre class="contents "><span class="cmd command">
sleep 100 &amp;
echo $! &gt; /cgroup1/child1/cgroup.procs
</span></pre></div>
<p class="para">
Other administration is done through files in the cgroup directories.  For
instance, to freeze all tasks in child1,
  </p>
<div class="screen"><pre class="contents "><span class="cmd command">
echo FROZEN &gt; /cgroup1/child1/freezer.state
</span></pre></div>
<p class="para">
A great deal of information about cgroups and its subsystems can be found
under the cgroups documentation directory in the kernel source tree (see
Resources).
  </p>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups-overview.html" title="Översikt">Föregående</a><a class="nextlinks-next" href="cgroups-delegation.html" title="Delegation">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
