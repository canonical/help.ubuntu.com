<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Växla mellan fönster</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord</a> › <a class="trail" href="shell-overview.html#apps" title="Program och fönster">Program och fönster</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord</a> › <a class="trail" href="shell-overview.html#apps" title="Program och fönster">Program och fönster</a> » <a class="trail" href="shell-windows.html" title="Fönster och arbetsytor">Fönster och arbetsytor</a> › <a class="trail" href="shell-windows.html#working-with-windows" title="Arbeta med fönster">Fönster</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Växla mellan fönster</span></h1></div>
<div class="region">
<div class="contents"></div>
<div id="launcher" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Från Startaren</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Visa <span class="gui">Programstartaren</span> genom att flytta din mus till din skärms övre vänstra hörn.</p></li>
<li class="steps"><p class="p">Öppna program har en liten vit triangulär pil till vänster. Klicka på ett öppet program för att växla till det.</p></li>
<li class="steps"><p class="p">Om ett öppet program har flera fönster öppna kommer det finnas många vita pilar till vänster. Klicka på programikonen en andra gång för att visa alla öppna fönster utzoomade. Klicka sedan på fönstret du vill växla till.</p></li>
</ol></div></div></div></div></div>
</div></div>
<div id="keyboard" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Från tangentbordet</span></h2></div>
<div class="region"><div class="contents">
<div class="list"><div class="inner"><div class="region"><ul class="list"><li class="list">
<p class="p">Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span> för att öppna <span class="gui">fönstervöxlaren</span>.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Släpp <span class="key"><kbd>Alt</kbd></span> för att välja nästa (markerade) fönster i växlaren.</p></li>
<li class="list">
<p class="p">Fortsätt annars hålla nere <span class="key"><kbd>Alt</kbd></span>-tangenten, och tryck <span class="key"><kbd>Tab</kbd></span> för att stega igenom listan över öppna fönster, eller <span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span> för att stega baklänges.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Fönster i fönsterväxlaren grupperas efter program. Miniatyrbilder av program med flera fönster dyker upp allt eftersom du klickar dig fram.</p></div></div></div></div>
</li>
<li class="list"><p class="p">Du kan också flytta mellan programikonerna i fönsterväxlaren med <span class="key"><kbd>→</kbd></span>- eller <span class="key"><kbd>←</kbd></span>-tangenterna eller välja en genom att klicka på den med musen.</p></li>
<li class="list">
<p class="p">Förhandsvisningar av program med ett enda fönster kan visas med <span class="key"><kbd>↓</kbd></span>-tangenten.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Bara fönster från den aktuella <span class="link"><a href="shell-workspaces.html" title="Vad är en arbetsyta, och vad har jag för nytta av den?">arbetsytan</a></span> kommer visas. För att visa fönster från alla arbetsytor, håll nere <span class="key"><kbd>Ctrl-</kbd></span> och <span class="key"><kbd>Alt-</kbd></span>tangenterna och tryck <span class="key"><kbd>Tab</kbd></span> eller <span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span>.</p></div></div></div></div>
</li>
</ul></div></div></div>
</li></ul></div></div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list"><li class="list">
<p class="p">Tryck <span class="keyseq"><span class="key"><kbd><span class="link"><a href="windows-key.html" title='Vad är "Superknappen"?'>Super</a></span></kbd></span>+<span class="key"><kbd>W</kbd></span></span> för att visa alla öppna fönster utzoomade.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list"><li class="list"><p class="p">Klicka på fönstret du vill växla till.</p></li></ul></div></div></div>
</li></ul></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="shell-windows.html#working-with-windows" title="Arbeta med fönster">Arbeta med fönster</a></li>
<li class="links "><a href="shell-overview.html#apps" title="Program och fönster">Program och fönster</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
