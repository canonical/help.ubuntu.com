�PNG

   IHDR      8   2�l1    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<  PLTE   ���������---������ttt$$$���bbb��������֦��ccc���QQQ���������������999���qqq���TTTJJJ���������%%%������������ddd���PPPKKK���)))���FFF���777888���;;;ooo>>>(((LLL������


�����Ө��������������aaa���mmm���'''���AAABBB���HHHhhh���vvvyyywww			   ��킂������������������ľ��ggg���SSSnnn___������,,,������&&&���RRRUUU������***��ɒ��[[[���������:::555������DDD��̑����»�����ppp���rrrEEE���CCC333���...~~~<<<���uuu���OOO}}}000��ݓ�����GGGIII4440q������7   bKGD�Cd��   tIME�	:��   caNv     X        QVz�  !IDATx����_Su��/_�/:��T`Ҝ���[�E�6��E�a8�bqGIRC-�]#b�����bg;g�m��8�����/|?�/������{�g         ���@�fkٺ�%:��)��(RŢH���= i�C-5���H�X��&��YZ�1O�k���-[�sz�+*eJeE9�x���U)�~_��ƣ�����PQ0��������\�ӫ}��ޝ������
i��s�����'P��UX�z���-k�c���(�i�(2�5I�\ֲwoKY��EM9��R�P;
]���u�]a٪7�˰�|TJ+�7��wt`5Z�'��f# �TI��QOls�8�Tg��g�<�ܡ�_X<����KZ+Ug���H��r����;��&#$_���#�����!��Z����c���v���9�z5���co�jz���mo��D@��:T�'��Q888�2���a��q��hsf_��8%�i��U$�D@��t�5c\��muF�+�ƵuC���
qN��w'�5�;`2�*�(�E�Q���mZ��ȍ��i�>�V��زT@.�U�z?U~Я��IqJ��*�ڳkpS΀��W���:��!�����W;�5뀌��������YJ���#����nrAV��GF]��q@}rD�mд����3�S=?�����	�0�j�K���1���p��C��X���r��Y"����������lガ$ ��z��	1�f�?�/\���rr.g�Ȝ&��hQj�Y�f5�|"1���Ns�>b�I/�*$���9G]oW��7`����=��_��I�o�u�+׵���w^�Y�(a<LM��Qd5� !e"o������<�y���g���?�Y��Q�T���{%BT_�����V�qϯ�	ˀA@lę�#���k��ب���_�܃`�����=��jrH��T�[2�dmZg�8Ԧ_r��)所 [[m���0J>        k�_ ,��    @@ ��    @@ ��    @@ �_�7Lg����Q   'tEXtCreation Time 2025-04-09T15:07:58-00:004�]   %tEXtdate:create 2025-04-09T15:07:58-00:00��x   %tEXtdate:modify 2025-04-09T15:07:58-00:00����   (tEXtdate:timestamp 2025-04-09T15:07:58-00:00���o   tEXtSoftware gnome-screenshot��>    IEND�B`�