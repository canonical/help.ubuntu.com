<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Why does my wireless network keep disconnecting?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-problem.html" title="Nätverksproblem">Nätverksproblem</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Why does my wireless network keep disconnecting?</span></h1></div>
<div class="region">
<div class="contents"><p class="p">You may find that you have been disconnected from a wireless network even though you wanted to stay connected. Your computer will normally try to reconnect to the network as soon as this happens (the network icon on the menu bar will pulse if it is trying to reconnect), but it can be annoying, especially if you were using the internet at the time.</p></div>
<div id="signal" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Weak wireless signal</span></h2></div>
<div class="region"><div class="contents">
<p class="p">A common reason for being disconnected from a wireless network is that you have low signal. Wireless networks have a limited range, so if you are too far away from the wireless base station you may not be able to get a strong enough signal to maintain a connection. Walls and other objects between you and the base station can also weaken the signal.</p>
<p class="p">The network icon on the menu bar displays how strong your wireless signal is. If the signal looks low, try moving closer to the wireless base station.</p>
</div></div>
</div></div>
<div id="network" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Network connection not being established properly</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Sometimes, when you connect to a wireless network, it may appear that you have successfully connected at first, but then you will be disconnected soon after. This normally happens because your computer was only partially successful in connecting to the network - it managed to establish a connection, but was unable to finalize the connection for some reason and so was disconnected.</p>
<p class="p">A possible reason for this is that you entered the wrong wireless passphrase, or that your computer was not allowed on the network (because the network requires a username to log in, for example).</p>
</div></div>
</div></div>
<div id="hardware" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Unreliable wireless hardware/drivers</span></h2></div>
<div class="region"><div class="contents"><p class="p">Some wireless network hardware can be a little unreliable. Wireless networks are complicated, so wireless cards and base stations occasionally run into minor problems and may drop connections. This is annoying, but it happens quite regularly with many devices. If you are disconnected from wireless connections from time to time, this may be the only reason. If it happens very regularly, you may want to consider getting some different hardware.</p></div></div>
</div></div>
<div id="busy" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Busy wireless networks</span></h2></div>
<div class="region"><div class="contents"><p class="p">Wireless networks in busy places (in universities and coffee shops, for example) often have many computers trying to connect to them at once. Sometimes these networks get too busy and may not be able to handle all of the computers that are trying to connect, so some of them get disconnected.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="net-problem.html" title="Nätverksproblem">Nätverksproblem</a><span class="desc"> — 
      <span class="link"><a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Troubleshooting wireless connections</a></span>,
      <span class="link"><a href="net-wireless-find.html" title="I can't see my wireless network in the list">finding your wifi network</a></span>…
        </span>
</li>
<li class="links ">
<a href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a><span class="desc"> — 
      <span class="link"><a href="net-wireless-connect.html" title="Connect to a wireless network">Connect to wifi</a></span>,
      <span class="link"><a href="net-wireless-hidden.html" title="Connect to a hidden wireless network">Hidden networks</a></span>,
      <span class="link"><a href="net-wireless-edit-connection.html" title="Redigera en trådlös anslutning">Edit connection settings</a></span>,
      <span class="link"><a href="net-wireless-disconnecting.html" title="Why does my wireless network keep disconnecting?">Disconnecting</a></span>…
    </span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless-connect.html" title="Connect to a wireless network">Connect to a wireless network</a><span class="desc"> — Get on the internet - wirelessly.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
