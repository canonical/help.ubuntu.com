<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Fönster och arbetsytor</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html.sv" title="Ditt skrivbord">Skrivbord</a> › <a class="trail" href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Fönster och arbetsytor</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Precis som andra skrivbord använder GNOME fönster för att visa dina körande program. Genom att använda både översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och <span class="em">snabbstartspanelen</span> kan du starta nya program och kontrollera aktiva fönster.</p>
<p class="p">Du kan också gruppera ihop dina program inom arbetsytor. Titta på hjälptexterna om fönster och arbetsytor nedan för att bättre förstår hur du använder dessa funktioner.</p>
</div>
<div id="working-with-windows" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Arbeta med fönster</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-windows-states.html.sv" title="Flytta och storleksändra fönster"><span class="title">Flytta och storleksändra fönster</span><span class="linkdiv-dash"> — </span><span class="desc">Ordna fönster på en arbetsyta för du ska kunna arbeta effektivare.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-windows-lost.html.sv" title="Hitta ett förlorat fönster"><span class="title">Hitta ett förlorat fönster</span><span class="linkdiv-dash"> — </span><span class="desc">Kontrollera översiktsvyn <span class="gui">Aktiviteter</span> eller andra arbetsytor.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-windows-maximize.html.sv" title="Maximera och avmaximera ett fönster"><span class="title">Maximera och avmaximera ett fönster</span><span class="linkdiv-dash"> — </span><span class="desc">Dubbelklicka på eller dra i en namnlist för att maximera eller återställa ett fönster.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-windows-tiled.html.sv" title="Placera fönster sida-vid-sida"><span class="title">Placera fönster sida-vid-sida</span><span class="linkdiv-dash"> — </span><span class="desc">Maximera två fönster sida-vid-sida.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-windows-switching.html.sv" title="Växla mellan fönster"><span class="title">Växla mellan fönster</span><span class="linkdiv-dash"> — </span><span class="desc">Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span>.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="working-with-workspaces" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Arbeta med arbetsytor</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-workspaces.html.sv" title="Vad är en arbetsyta, och hur hjälper den mig?"><span class="title">Vad är en arbetsyta, och hur hjälper den mig?</span><span class="linkdiv-dash"> — </span><span class="desc">Arbetsytor är ett sätta gruppera fönster på ditt skrivbord.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-workspaces-movewindow.html.sv" title="Flytta ett fönster till en annan arbetsyta"><span class="title">Flytta ett fönster till en annan arbetsyta</span><span class="linkdiv-dash"> — </span><span class="desc">Gå till översiktsvyn <span class="gui">Aktiviteter</span> och dra fönstret till en annan arbetsyta.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="shell-workspaces-switch.html.sv" title="Växla mellan arbetsytor"><span class="title">Växla mellan arbetsytor</span><span class="linkdiv-dash"> — </span><span class="desc">Använd arbetsyteväxlaren.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
