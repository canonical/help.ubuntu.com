<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Komma igång</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 19.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Komma igång</span></h1></div>
<div class="region"><div class="contents">
<div class="ui-tile ">
<a href="figures/gnome-launching-applications.webm" class="ui-overlay"><span class="ui-tile-img" style="width: 235px; height: 145px;"><img src="gs-thumb-launching-apps.svg" width="235" height="145"></span><span class="ui-tile-text" style="max-width: 235px;"><span class="desc center">Starta program</span></span></a><div class="ui-overlay"><div class="inner">
<a href="#" class="ui-overlay-close" title="Stäng">⨯</a><div class="contents"><div class="media media-video"><div class="inner">
<video src="figures/gnome-launching-applications.webm" preload="auto" controls="controls" class="media media-block" height="394" width="700" data-play-label="Spela upp" data-pause-label="Paus"></video><div class="media-ttml">
<div class="media-ttml-node media-ttml-div" data-ttml-begin="1" data-ttml-end="5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="1" data-ttml-end="5">Starta program</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="5" data-ttml-end="7.5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="5" data-ttml-end="7.5">Flytta din musmarkör till <span class="gui">Aktivitetshörnet</span> längst upp till vänster på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="7.5" data-ttml-end="9.5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="7.5" data-ttml-end="9.5">Klicka på ikonen <span class="gui">Visa program</span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="9.5" data-ttml-end="11"><div class="media-ttml-node media-ttml-p" data-ttml-begin="9.5" data-ttml-end="11">Klicka på programmet som du vill köra, till exempel, Hjälp.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="12" data-ttml-end="21"><div class="media-ttml-node media-ttml-p" data-ttml-begin="12" data-ttml-end="21">Alternativt, använd tangentbordet för att öppna <span class="gui">Aktivitetsöversikt</span> genom att trycka på <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="22" data-ttml-end="29"><div class="media-ttml-node media-ttml-p" data-ttml-begin="22" data-ttml-end="29">Börja skriva namnet på det program du vill starta.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="30" data-ttml-end="33"><div class="media-ttml-node media-ttml-p" data-ttml-begin="30" data-ttml-end="33">Tryck på <span class="key"><kbd>Retur</kbd></span> för att starta programmet.</div></div>
</div>
</div></div></div>
</div></div>
</div>
<div class="ui-tile ">
<a href="figures/gnome-task-switching.webm" class="ui-overlay"><span class="ui-tile-img" style="width: 235px; height: 145px;"><img src="gs-thumb-task-switching.svg" width="235" height="145"></span><span class="ui-tile-text" style="max-width: 235px;"><span class="desc center">Växla uppgifter</span></span></a><div class="ui-overlay"><div class="inner">
<a href="#" class="ui-overlay-close" title="Stäng">⨯</a><div class="contents"><div class="media media-video"><div class="inner">
<video src="figures/gnome-task-switching.webm" preload="auto" controls="controls" class="media media-block" height="394" width="700" data-play-label="Spela upp" data-pause-label="Paus"></video><div class="media-ttml">
<div class="media-ttml-node media-ttml-div" data-ttml-begin="1" data-ttml-end="5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="1" data-ttml-end="5">Växlar uppgifter</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="5" data-ttml-end="8"><div class="media-ttml-node media-ttml-p" data-ttml-begin="5" data-ttml-end="8">Flytta din musmarkör till <span class="gui">Aktivitetshörnet</span> längst upp till vänster på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="9" data-ttml-end="12"><div class="media-ttml-node media-ttml-p" data-ttml-begin="9" data-ttml-end="12">Klicka på ett fönster för att byta till den uppgiften.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="12" data-ttml-end="14"><div class="media-ttml-node media-ttml-p" data-ttml-begin="12" data-ttml-end="14">För att maximera ett fönster längs skärmens vänstra sida, fånga fönstrets namnlist och dra det åt vänster.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="14" data-ttml-end="16"><div class="media-ttml-node media-ttml-p" data-ttml-begin="14" data-ttml-end="16">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="16" data-ttml-end="0"><div class="media-ttml-node media-ttml-p" data-ttml-begin="16" data-ttml-end="0">För att maximera ett fönster längs den högra sidan, fånga fönstrets namnlist och dra det åt höger.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="18" data-ttml-end="20"><div class="media-ttml-node media-ttml-p" data-ttml-begin="18" data-ttml-end="20">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="23" data-ttml-end="27"><div class="media-ttml-node media-ttml-p" data-ttml-begin="23" data-ttml-end="27">Tryck <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>+<span class="key"><kbd> Tabb</kbd></span></span> för att visa <span class="gui">fönsterväxlaren</span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="27" data-ttml-end="29"><div class="media-ttml-node media-ttml-p" data-ttml-begin="27" data-ttml-end="29">Släpp <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> för att välja nästa markerade fönster.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="29" data-ttml-end="32"><div class="media-ttml-node media-ttml-p" data-ttml-begin="29" data-ttml-end="32">För att bläddra igenom listan av öppna fönster, släpp inte <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> utan håll den nertryckt och tryck på <span class="key"><kbd>Tabb</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="35" data-ttml-end="37"><div class="media-ttml-node media-ttml-p" data-ttml-begin="35" data-ttml-end="37">Tryck på <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super </kbd></a></span> för att visa <span class="gui">Aktivitetsöversikt</span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="37" data-ttml-end="40"><div class="media-ttml-node media-ttml-p" data-ttml-begin="37" data-ttml-end="40">Börja skriv in namnet på det program du vill växla till.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="40" data-ttml-end="43"><div class="media-ttml-node media-ttml-p" data-ttml-begin="40" data-ttml-end="43">När programmet visas som det första resultatet, tryck på <span class="key"><kbd>Retur</kbd></span> för att växla till det.</div></div>
</div>
</div></div></div>
</div></div>
</div>
<div class="ui-tile ">
<a href="figures/gnome-windows-and-workspaces.webm" class="ui-overlay"><span class="ui-tile-img" style="width: 235px; height: 145px;"><img src="gs-thumb-windows-and-workspaces.svg" width="235" height="145"></span><span class="ui-tile-text" style="max-width: 235px;"><span class="desc center">Använda fönster och arbetsytor</span></span></a><div class="ui-overlay"><div class="inner">
<a href="#" class="ui-overlay-close" title="Stäng">⨯</a><div class="contents"><div class="media media-video"><div class="inner">
<video src="figures/gnome-windows-and-workspaces.webm" preload="auto" controls="controls" class="media media-block" height="394" width="700" data-play-label="Spela upp" data-pause-label="Paus"></video><div class="media-ttml">
<div class="media-ttml-node media-ttml-div" data-ttml-begin="1" data-ttml-end="5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="1" data-ttml-end="5">Fönster och arbetsytor</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="6" data-ttml-end="10"><div class="media-ttml-node media-ttml-p" data-ttml-begin="6" data-ttml-end="10">För att maximera ett fönster, fånga fönstrets namnlist och dra det till toppen på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="10" data-ttml-end="13"><div class="media-ttml-node media-ttml-p" data-ttml-begin="10" data-ttml-end="13">När skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="14" data-ttml-end="20"><div class="media-ttml-node media-ttml-p" data-ttml-begin="14" data-ttml-end="20">För att avmaximera ett fönster, fånga fönstrets namnlist och dra det bort ifrån kanterna på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="25" data-ttml-end="29"><div class="media-ttml-node media-ttml-p" data-ttml-begin="25" data-ttml-end="29">Du kan också klicka på namnlisten för att dra bort fönstret och avmaximera det.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="34" data-ttml-end="38"><div class="media-ttml-node media-ttml-p" data-ttml-begin="34" data-ttml-end="38">För att maximera ett fönster längs skärmens vänstra sida, fånga fönstrets namnlist och dra det åt vänster.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="38" data-ttml-end="40"><div class="media-ttml-node media-ttml-p" data-ttml-begin="38" data-ttml-end="40">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="41" data-ttml-end="44"><div class="media-ttml-node media-ttml-p" data-ttml-begin="41" data-ttml-end="44">För att maximera ett fönster längs skärmens högra sida, fånga fönstrets namnlist och dra det åt höger.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="44" data-ttml-end="48"><div class="media-ttml-node media-ttml-p" data-ttml-begin="44" data-ttml-end="48">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="54" data-ttml-end="60"><div class="media-ttml-node media-ttml-p" data-ttml-begin="54" data-ttml-end="60">För att maximera ett fönster med tangentbordet, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>↑</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="61" data-ttml-end="66"><div class="media-ttml-node media-ttml-p" data-ttml-begin="61" data-ttml-end="66">För att återställa fönstret till dess avmaximerade storlek, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>↓</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="66" data-ttml-end="73"><div class="media-ttml-node media-ttml-p" data-ttml-begin="66" data-ttml-end="73">För att maximera ett fönster längs den högra sidan på skärmen, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>→</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="76" data-ttml-end="82"><div class="media-ttml-node media-ttml-p" data-ttml-begin="76" data-ttml-end="82">För att maximera ett fönster längs den vänstra sidan på skärmen, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>←</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="83" data-ttml-end="89"><div class="media-ttml-node media-ttml-p" data-ttml-begin="83" data-ttml-end="89">För att flytta till en arbetsyta som är under den nuvarande arbetsytan, tryck på <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super </kbd></a></span>+<span class="key"><kbd>Page Down</kbd></span></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="90" data-ttml-end="97"><div class="media-ttml-node media-ttml-p" data-ttml-begin="90" data-ttml-end="97">För att flytta till en arbetsyta som är ovanför den nuvarande arbetsytan, tryck på <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super </kbd></a></span>+<span class="key"><kbd>Page Up</kbd></span></span>.</div></div>
</div>
</div></div></div>
</div></div>
</div>
<div class="links topiclinks"><div class="inner">
<div class="title title-links title-heading"><h2><span class="title">Vanliga uppgifter</span></h2></div>
<div class="region">
<div class="links-grid "><div class="links-grid-link"><a href="gs-connect-online-accounts.html.sv" title="Ansluta till nätkonton">Ansluta till nätkonton</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-use-system-search.html.sv" title="Använd systemsökning">Använd systemsökning</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-use-windows-workspaces.html.sv" title="Använda fönster och arbetsytor">Använda fönster och arbetsytor</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-browse-web.html.sv" title="Surfa på nätet">Surfa på nätet</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-change-wallpaper.html.sv" title="Ändra bakgrund">Ändra bakgrund</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-change-date-time-timezone.html.sv" title="Ändra datum, tid och tidszon">Ändra datum, tid och tidszon</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-get-online.html.sv" title="Ansluta till nätet">Ansluta till nätet</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-launch-applications.html.sv" title="Starta program">Starta program</a></div></div>
<div class="links-grid "><div class="links-grid-link"><a href="gs-switch-tasks.html.sv" title="Växla uppgifter">Växla uppgifter</a></div></div>
</div>
</div></div>
<div class="links guidelinks"><div class="inner">
<div class="title title-links"><h2><span class="title"></span></h2></div>
<div class="region"><ul class="links-heading"><li class="links "><div class="links-heading"><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></div></li></ul></div>
</div></div>
</div></div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
