<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Hantera program &amp; inställningar via menypanelen</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Hantera program &amp; inställningar via menypanelen</span></h1></div>
<div class="region">
<div class="contents"><p class="p">The <span class="gui">menu bar</span> is the dark strip on the top of your screen.
    It contains the window management buttons, the app menus, and the status menus.</p></div>
<div id="window-management" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Window management buttons</span></h2></div>
<div class="region">
<div class="contents"><p class="p">The <span class="gui">window management buttons</span> are on the top left corner of windows. When
    maximized, the buttons are in the top left of the screen. Click the buttons to
    close, minimize, maximize or restore windows.</p></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="shell-windows-states.html" title="Window operations">Window operations</a><span class="desc"> — Restore, resize, arrange and hide.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="app-menus" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Programmenyer</span></h2></div>
<div class="region"><div class="contents">
<p class="p">The <span class="gui">app menus</span> are by default located to the right of the window management buttons.
    Unity hides the app menus and the window management buttons unless you move your
    mouse pointer to the top left of the screen or press <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F10</kbd></span></span>.
    This feature enables you to see more of your content at once, which is
    especially valuable on small screens like netbooks.
  </p>
<p class="p">If you want, you can change the default behavior, and have your menus attached
    to the window title bar of respective application instead of the menu bar.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ikonen längst till höger i menyraden och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">In the Personal section, click <span class="gui">Appearance</span> and choose the
        <span class="gui">Behavior</span> tab.</p></li>
<li class="steps"><p class="p">Under <span class="gui">Show the menus for a window</span>, select <span class="gui">In the window's title bar</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="status-menus" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Statusmenyer</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Ubuntu has several different <span class="gui">status menus</span> (sometimes referred to as
    <span class="gui">indicators</span>) on the right side of the menu bar.
    The status menus are a convenient place where you can check and modify the
    state of your computer and applications.</p>
<div class="list ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-list"><h3><span class="title">List of status menus and what they do</span></h3></div>
<div class="region"><ul class="list">
<li class="list">
<p class="p"><span class="em">Network menu</span> <span class="media"><span class="media media-image"><img src="img/network-offline.svg" class="media media-inline" alt="Offline network icon"></span></span></p>
<p class="p">Connect to <span class="link"><a href="net-wired-connect.html" title="Connect to a wired (Ethernet) network">wired</a></span>, <span class="link"><a href="net-wireless-connect.html" title="Connect to a wireless network">wireless</a></span>,
        <span class="link"><a href="net-mobile.html" title="Connect to mobile broadband">mobile</a></span>, and <span class="link"><a href="net-vpn-connect.html" title="Connect to a VPN">VPN</a></span> networks.</p>
</li>
<li class="list">
<p class="p"><span class="em">Input source menu</span> <span class="media"><span class="media media-image"><img src="img/indicator-keyboard-En.svg" class="media media-inline" alt="Input source icon"></span></span></p>
<p class="p">Select keyboard layout/input source, <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">configure input sources</a></span>.</p>
</li>
<li class="list">
<p class="p"><span class="em">Bluetooth menu</span> <span class="media"><span class="media media-image"><img src="img/bluetooth-active.svg" class="media media-inline" alt="Bluetooth icon"></span></span></p>
<p class="p">Send or receive files by <span class="link"><a href="bluetooth.html" title="Bluetooth">Bluetooth</a></span>. This menu
        is hidden if a supported Bluetooth device isn't detected.</p>
</li>
<li class="list">
<p class="p"><span class="em">Messaging menu</span> <span class="media"><span class="media media-image"><img src="img/indicator-messages.svg" class="media media-inline" alt="Message icon"></span></span></p>
<p class="p">Easily launch and receive incoming notifications from messaging applications
         including email, social networking, and Internet chat.</p>
</li>
<li class="list">
<p class="p"><span class="em">Battery menu</span> <span class="media"><span class="media media-image"><img src="img/battery-100.svg" class="media media-inline" alt="Battery icon"></span></span></p>
<p class="p">Check your laptop battery's charging status. This menu is
       hidden if a battery isn't detected.</p>
</li>
<li class="list">
<p class="p"><span class="em">Sound menu</span> <span class="media"><span class="media media-image"><img src="img/audio-volume-high-panel.svg" class="media media-inline" alt="Volume icon"></span></span></p>
<p class="p">Set the <span class="link"><a href="sound-volume.html" title="Change the sound volume">volume</a></span>, configure sound <span class="link"><a href="media.html" title="Ljud, video och bilder">settings</a></span>,
        and control media players like <span class="app">Rhythmbox</span>.</p>
</li>
<li class="list">
<p class="p"><span class="em">Clock</span></p>
<p class="p">Access the current time and date. Appointments from your
        <span class="link"><a href="clock-calendar.html" title="Kalendermöten">Evolution calendar</a></span> can also display here.</p>
</li>
<li class="list">
<p class="p"><span class="em">System menu</span> <span class="media"><span class="media media-image"><img src="img/system-devices-panel.svg" class="media media-inline" alt="Power cog icon"></span></span></p>
<p class="p">Access details about your computer, this help guide, and <span class="link"><a href="prefs.html" title="Inställningar för användare och system">system settings</a></span>.
        Switch users, lock screen, log out, suspend, restart or shutdown your computer.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Some of the icons used by the indicator menus change according to the status of the application.</p></div></div></div></div>
<p class="p">Other programs such as <span class="app">Tomboy</span> or <span class="app">Transmission</span> can also add indicator menus to the panel.</p>
</li>
</ul></div>
</div>
</div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
