<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Referenser</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="package-management.html" title="Pakethantering">Pakethantering</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="configuration.html" title="Konfiguration">Föregående</a><a class="nextlinks-next" href="networking.html" title="Nätverk">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Referenser</h1></div>
<div class="region"><div class="contents">
<p class="para">De mesta av materialet som ingår i detta kapitel finns i <span class="app application">man</span>-sidorna, många av dessa är tillgängliga på nätet.</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
        <p class="para">
        The <a href="https://help.ubuntu.com/community/InstallingSoftware" class="ulink" title="https://help.ubuntu.com/community/InstallingSoftware">InstallingSoftware</a> Ubuntu wiki page has more information.
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        For more <span class="app application">dpkg</span> details see the 
        <a href="http://manpages.ubuntu.com/manpages/trusty/en/man1/dpkg.1.html" class="ulink" title="http://manpages.ubuntu.com/manpages/trusty/en/man1/dpkg.1.html">dpkg man page</a>.
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        The <a href="http://www.debian.org/doc/manuals/apt-howto/" class="ulink" title="http://www.debian.org/doc/manuals/apt-howto/">APT HOWTO</a> and 
        <a href="http://manpages.ubuntu.com/manpages/trusty/en/man8/apt-get.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/trusty/en/man8/apt-get.8.html">apt-get man page</a>
        contain useful information regarding <span class="app application">apt-get</span> usage.
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">
        See the <a href="http://manpages.ubuntu.com/manpages/trusty/man8/aptitude.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/trusty/man8/aptitude.8.html">aptitude man page</a> 
        for more <span class="app application">aptitude</span> options.
        </p>
      </li>
<li class="list itemizedlist">
        <p class="para">Sidan <a href="https://help.ubuntu.com/community/Repositories/Ubuntu" class="ulink" title="https://help.ubuntu.com/community/Repositories/Ubuntu">Adding Repositories HOWTO (Ubuntu Wiki)</a> innehåller mer detaljer om att lägga till förråd.</p>
      </li>
</ul></div>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="configuration.html" title="Konfiguration">Föregående</a><a class="nextlinks-next" href="networking.html" title="Nätverk">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
