<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Välj ett säkert lösenord</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="user-accounts.html.sv" title="Användarkonton">Användare</a> › <a class="trail" href="user-accounts.html.sv#passwords" title="Lösenord">Lösenord</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Välj ett säkert lösenord</span></h1></div>
<div class="region">
<div class="contents">
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">Gör dina lösenord enkla nog för att själv komma ihåg dem, men svåra för andra (inklusive datorprogram) att gissa.</p></div></div></div></div>
<p class="p">Att välja ett bra lösenord kommer att hjälpa till att hålla din dator säker. Om lösenordet är lätt att gissa kan någon komma på det och få tillgång till din personliga information.</p>
<p class="p">Personer kan till och med använda datorer för att systematiskt försöka gissa ditt lösenord, så även ett som skulle vara svårt för en människa att gissa kan vara extremt enkelt för ett datorprogram att knäcka. Här kommer några tips om hur du väljer ett bra lösenord:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list">
<p class="p">Använd en blandning av stora och små bokstäver, siffror symboler och mellanslag i lösenordet. Detta gör det svårare att gissa; det finns fler symboler att välja mellan vilket innebär fler möjliga lösenord som någon måste kontrollera när de försöka gissa ditt.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Ett bra sätt för att välja ett lösenord är att ta den första bokstaven i varje ord i en fras som du kan komma ihåg. Frasen kan vara namnet på en film, en bok, en låt eller ett album. Till exempel skulle ”Flatland: A Romance of Many Dimensions” bli F:ARoMD eller faromd eller f: aromd.</p></div></div></div></div>
</li>
<li class="list"><p class="p">Gör dina lösenord så långa som möjligt. Ju fler tecken det innehåller, desto längre bör det ta för en person eller dator att gissa det.</p></li>
<li class="list"><p class="p">Använd inte några ord som dyker upp i ett standarduppslagsverk på något språk. Lösenordsknäckare kommer att försöka med dessa först. Det vanligaste lösenordet är ”password” — personer kan gissa lösenord som detta väldigt snabbt!</p></li>
<li class="list"><p class="p">Använd inte någon personlig information så som datum, registreringsnummer eller familjemedlemmars namn.</p></li>
<li class="list"><p class="p">Använd inte några substantiv.</p></li>
<li class="list">
<p class="p">Välj ett lösenord som kan skriva snabbt, för att minska chanserna att någon kan lista ut vad du skrivit om de råkar se dig.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Skriv aldrig ner dina lösenord någonstans. De kan hittas lätt!</p></div></div></div></div>
</li>
<li class="list"><p class="p">Använd olika lösenord för olika saker.</p></li>
<li class="list">
<p class="p">Använd olika lösenord för olika konton.</p>
<p class="p">Om du använder samma lösenord för alla dina konton, kan den som listar ut det omedelbart få tillgång till alla dina konton.</p>
<p class="p">Det kan dock vara svårt att komma ihåg många lösenord. Även om det inte är lika säkert som att välja olika lösenord för allting så kan det vara lättare att använda samma för saker som inte spelar någon roll (som webbplatser), och olika för viktiga saker (som din internetbank och din e-post).</p>
</li>
<li class="list"><p class="p">Byt dina lösenord regelbundet.</p></li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="user-accounts.html.sv#passwords" title="Lösenord">Lösenord</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="user-changepassword.html.sv" title="Välj ditt lösenord">Välj ditt lösenord</a><span class="desc"> — Håll ditt konto säkert genom att ändra ditt lösenord ofta i dina kontoinställningar.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
