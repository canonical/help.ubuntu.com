<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="500" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-search-settings.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17453" ns4:href="#linearGradient5716" ns1:collect="always"/>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17455" ns4:href="#linearGradient5716" ns1:collect="always"/>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2-0">
      <ns0:stop id="stop3964-5-0-1-9-6-6-34" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6-4" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7-0"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3-6" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath15654">
      <ns0:path ns2:type="arc" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.99999994;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="path15656" ns2:cx="180.375" ns2:cy="183.625" ns2:rx="20.875" ns2:ry="20.875" d="m 201.25,183.625 a 20.875,20.875 0 1 1 -41.75,0 A 20.875,20.875 0 1 1 201.25,183.625 Z" transform="translate(253.75,41.5)"/>
    </ns0:clipPath>
    <ns0:filter style="color-interpolation-filters:sRGB" height="1.1308649" id="filter5601" width="1.2058235" x="-0.10291173" y="-0.065432459" ns1:collect="always">
      <ns0:feGaussianBlur id="feGaussianBlur5603" stdDeviation="0.610872" ns1:collect="always"/>
    </ns0:filter>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5176" gradientUnits="userSpaceOnUse" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath5304">
      <ns0:rect ry="0.1367164" rx="0.26726839" y="638.97058" x="606.59344" height="136.72638" width="141.10645" id="rect5306" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.50848383;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath987">
      <ns0:circle r="60" cy="236" cx="63.999996" id="circle989" style="display:inline;opacity:1;fill:#3584e4;fill-opacity:1;stroke:none;stroke-width:4.28571415;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath987-2">
      <ns0:circle r="60" cy="236" cx="63.999996" id="circle989-0" style="display:inline;opacity:1;fill:#3584e4;fill-opacity:1;stroke:none;stroke-width:4.28571415;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="442.64988" ns1:cy="142.83514" ns1:document-units="px" ns1:current-layer="g4890" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="2560" ns1:window-height="1376" ns1:window-x="0" ns1:window-y="27" ns1:window-maximized="1" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="656" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-540)">
    <ns0:g style="display:inline" id="g4890" transform="matrix(2.6833333,0,0,2.6833333,-1275.5101,-1072.8539)">
      <ns0:path style="display:inline;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-opacity:1" d="m 506.43234,611.75299 h 258.32299 c 2.21601,0 4,1.784 4,4 v 161.2298 h -4 -258.32299 -4 v -161.2298 c 0,-2.216 1.784,-4 4,-4 z" id="path5430-2" ns1:connector-curvature="0" ns2:nodetypes="sssccccss"/>
      <ns0:path ns1:connector-curvature="0" id="path5361-7" d="M 502.98343,630.36169 H 768.47408" style="display:inline;fill:none;stroke:#000000;stroke-width:1.01455009;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:nodetypes="cc"/>
      <ns0:path style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.3358984;marker:none;enable-background:new" id="path5375-0" d="m 756.48074,617.84776 h 0.74998 c 0.008,-9e-5 0.0156,-3.5e-4 0.0234,0 0.19121,0.008 0.38239,0.0964 0.51561,0.23437 l 1.71089,1.71088 1.73432,-1.71088 c 0.19921,-0.17287 0.335,-0.22912 0.51561,-0.23437 h 0.74998 v 0.74998 c 0,0.21484 -0.0258,0.41297 -0.1875,0.56248 l -1.71088,1.71089 1.68745,1.68745 c 0.14113,0.14112 0.21092,0.34008 0.21093,0.53905 v 0.74997 h -0.74998 c -0.19897,0 -0.39793,-0.0698 -0.53905,-0.21093 l -1.71088,-1.71089 -1.71089,1.71089 c -0.14112,0.14114 -0.34009,0.21093 -0.53905,0.21093 h -0.74998 v -0.74997 c 0,-0.19897 0.0698,-0.39793 0.21094,-0.53905 l 1.71088,-1.68745 -1.71088,-1.71089 c -0.15806,-0.14597 -0.22737,-0.35193 -0.21094,-0.56248 z" ns1:connector-curvature="0" ns2:nodetypes="ccccccccscccccscccscsccccc"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:12px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1" x="669.13416" y="622.67841" id="text12012-9"><ns0:tspan ns2:role="line" id="tspan12014-3" x="669.13416" y="622.67841" style="font-size:5.21739101px;line-height:1.25;stroke-width:1">Sök</ns0:tspan></ns0:text>
      <ns0:rect width="5.9627328" height="5.9627328" x="-514.0741" y="617.82538" id="rect10837-5-8-1-6" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.3726708;marker:none;enable-background:new" transform="scale(-1,1)"/>
      <ns0:path d="m 512.58846,618.5707 h -0.37267 c -0.004,-4e-5 -0.008,-1.7e-4 -0.0117,0 -0.095,0.004 -0.19001,0.0479 -0.25621,0.11646 l -2.34696,2.13121 2.34698,2.13121 c 0.0701,0.0701 0.16899,0.10482 0.26786,0.10482 h 0.37267 v -0.37267 c 0,-0.0989 -0.0347,-0.19774 -0.10481,-0.26786 l -1.79962,-1.5955 1.79962,-1.59549 c 0.0785,-0.0725 0.11297,-0.17488 0.10481,-0.27951 z" ns1:connector-curvature="0" id="path10839-9-9-5-0" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.66381985;marker:none;enable-background:new" ns2:nodetypes="ccsccccccccccc"/>
      <ns0:rect style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.3726708;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" id="rect15386-6" width="11.925466" height="11.925466" x="505.35669" y="615.02728" rx="1.4906832" ry="1.4906832"/>
      <ns0:text id="text946" y="622.67841" x="541.68079" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:12px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1" xml:space="preserve"><ns0:tspan style="font-size:5.21739101px;line-height:1.25;stroke-width:1" y="622.67841" x="541.68079" id="tspan944" ns2:role="line">Inställningar</ns0:tspan></ns0:text>
      <ns0:rect transform="scale(-1,1)" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.3726708;marker:none;enable-background:new" id="rect948" y="617.82538" x="-575.56482" height="5.9627328" width="5.9627328"/>
      <ns0:rect ry="1.4906832" rx="1.4906832" y="615.02728" x="566.84741" height="11.925466" width="11.925466" id="rect952" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.3726708;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate"/>
      <ns0:g ns1:label="open-menu" id="g7352" transform="matrix(0.37267081,0,0,0.37267081,562.5214,515.34088)" style="display:inline;enable-background:new">
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" id="rect7354" width="16" height="16" x="20" y="276"/>
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7356" width="9.9996014" height="2.0002136" x="23.000198" y="278.99979"/>
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7358" width="9.9996014" height="2.0002136" x="23.000198" y="282.99979"/>
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7360" width="9.9996014" height="2.0002136" x="23.000198" y="286.99979"/>
      </ns0:g>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7822" width="79.006218" height="17.142857" x="502.92303" y="646.15674"/>
      <ns0:text id="text7826" y="656.21881" x="522.14331" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:12px;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:1" xml:space="preserve"><ns0:tspan style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.21739101px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;text-anchor:start;fill:#ffffff;stroke-width:1" y="656.21881" x="522.14331" id="tspan7824" ns2:role="line">Sök</ns0:tspan></ns0:text>
      <ns0:path style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" d="M 582.12691,611.30064 V 776.21886" id="path7828" ns1:connector-curvature="0"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7830" width="17.888199" height="3.3540373" x="521.92926" y="636.83997"/>
      <ns0:rect y="670.38031" x="521.92926" height="3.3540373" width="27.577641" id="rect7832" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7834" width="17.888199" height="3.3540373" x="521.92926" y="685.28717"/>
      <ns0:rect y="685.28717" x="544.28955" height="3.3540373" width="28.695652" id="rect7836" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="path7840" cx="511.71103" cy="638.71655" r="4.2555118"/>
      <ns0:circle r="4.2555118" cy="672.62958" cx="511.71103" id="circle7842" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle7844" cx="511.71103" cy="686.79108" r="4.2555118"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:7.45341635;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal" id="rect1222" width="2.6351805" height="45.325108" x="762.85754" y="634.08838" rx="1.3175902" ry="1.3175902"/>
      <ns0:rect width="5.9627328" height="5.9627328" x="509.25842" y="651.00146" id="rect3664" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.66372675;marker:none;enable-background:new"/>
      <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect3923-2" width="19.803892" height="10.92049" x="729.96857" y="615.98438" rx="5.4602423" ry="5.4602423"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="path915" cx="743.92047" cy="621.44116" r="4.4139271"/>
      <ns0:rect style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.50848383;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" id="rect12010-7" width="141.10643" height="137.72638" x="606.59344" y="638.97058" rx="0.26726839" ry="0.1367164"/>
      <ns0:g id="g5300" clip-path="url(#clipPath5304)">
        <ns0:rect ry="5.4602423" rx="5.4602423" y="646.65924" x="720.35028" height="10.92049" width="19.803892" id="rect3923-2-2" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
        <ns0:circle r="4.4139271" cy="652.11603" cx="734.30219" id="path915-5" style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect y="650.25616" x="634.84851" height="4.0993791" width="51.428574" id="rect5223" style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect5225" width="19.803892" height="10.92049" x="720.35028" y="661.5661" rx="5.4602423" ry="5.4602423"/>
        <ns0:circle style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5227" cx="734.30219" cy="667.02289" r="4.4139271"/>
        <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect5229" width="51.428574" height="4.0993791" x="634.84851" y="665.16302"/>
        <ns0:rect ry="5.4602423" rx="5.4602423" y="676.47296" x="720.35028" height="10.92049" width="19.803892" id="rect5231" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
        <ns0:circle r="4.4139271" cy="681.92975" cx="734.30219" id="circle5233" style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect y="680.06989" x="634.84851" height="4.0993791" width="51.428574" id="rect5235" style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect5237" width="19.803892" height="10.92049" x="720.35028" y="691.37982" rx="5.4602423" ry="5.4602423"/>
        <ns0:circle style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5239" cx="734.30219" cy="696.83661" r="4.4139271"/>
        <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect5241" width="51.428574" height="4.0993791" x="634.84851" y="694.97675"/>
        <ns0:rect ry="5.4602423" rx="5.4602423" y="706.28668" x="720.35028" height="10.92049" width="19.803892" id="rect5243" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
        <ns0:circle r="4.4139271" cy="711.74347" cx="734.30219" id="circle5245" style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect y="709.88361" x="634.84851" height="4.0993791" width="51.428574" id="rect5247" style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect5249" width="19.803892" height="10.92049" x="720.35028" y="721.19354" rx="5.4602423" ry="5.4602423"/>
        <ns0:circle style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5251" cx="734.30219" cy="726.65033" r="4.4139271"/>
        <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect5253" width="51.428574" height="4.0993791" x="634.84851" y="724.79047"/>
        <ns0:rect ry="5.4602423" rx="5.4602423" y="736.1004" x="720.35028" height="10.92049" width="19.803892" id="rect5255" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
        <ns0:circle r="4.4139271" cy="741.55719" cx="734.30219" id="circle5257" style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect y="739.69733" x="634.84851" height="4.0993791" width="51.428574" id="rect5259" style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect style="display:inline;fill:#deddda;fill-opacity:1;stroke:none;stroke-width:0.3726708" id="rect5261" width="19.803892" height="10.92049" x="720.35028" y="751.00726" rx="5.4602423" ry="5.4602423"/>
        <ns0:circle style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5263" cx="726.47607" cy="756.46405" r="4.4139271"/>
        <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect5265" width="51.428574" height="4.0993791" x="634.84851" y="754.60419"/>
        <ns0:rect ry="5.4602423" rx="5.4602423" y="765.91412" x="720.35028" height="10.92049" width="19.803892" id="rect5267" style="display:inline;fill:#deddda;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
        <ns0:circle r="4.4139271" cy="771.37091" cx="726.47607" id="circle5269" style="display:inline;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:rect y="769.51105" x="634.84851" height="4.0993791" width="51.428574" id="rect5271" style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:circle r="5.4913659" cy="711.74695" cx="622.92303" id="circle5329" style="display:inline;opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:circle style="display:inline;opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5331" cx="622.92303" cy="726.65381" r="5.4913659"/>
        <ns0:circle r="5.4913659" cy="741.56067" cx="622.92303" id="circle5333" style="display:inline;opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:circle style="display:inline;opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5335" cx="622.92303" cy="756.46753" r="5.4913659"/>
        <ns0:circle r="5.4913659" cy="771.37439" cx="622.92303" id="circle5337" style="display:inline;opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:g style="display:inline" id="g6180" transform="matrix(0.0931677,0,0,0.0931677,661.29603,605.68642)">
          <ns0:g style="display:inline;stroke-width:0.93333334;enable-background:new" transform="matrix(0.26785714,0,0,0.26785714,-482.48304,489.73394)" id="g912-6">
            <ns0:circle r="224" cy="43.999989" cx="256" id="circle1036" style="display:inline;opacity:1;fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:14.9333334;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
          </ns0:g>
          <ns0:path ns2:nodetypes="ccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccc" ns1:connector-curvature="0" id="path991" d="m 38,176 v 4 l 10,8 v 8 l 8,8 h 4 v -4 l 6,-6 v -4 l 4,-4 v -10 z m -4,16 H 4 c 0,0 0.5090211,40.4419 0,40 l 20,18 v -6 l -4,-4 6,-6 h 4 l 4,4 0.12494,-8.4018 L 40,224 h 4 v -4 l 4,-4 v -6 L 43.727619,206.12499 34,206 v 8 h -4 l -4,-4 v -4 l 6,-6 h 6 v -4 z m 60,2 -6,6 v 4 h 6 v -2.14287 h 4 v 4.26786 L 96,208 H 86 v 4 h -4 v 6 h -8 v 8 h 10 v -4 h 8 v 2 l 4,4 h 2 v -2 l -2,-2 v -2 h 4 l 6,6 h 6 v 2 l -2,2 h -4 l 18,18 V 194 H 96 Z m 12,38 H 94 l -2,-2 H 78 l -8,8 v 8 l 8,8 h 6 l 4,4 v 2 l 2,2 v 12 l 14,14 h 8 v -30 l 4,-4 v -8 l -10,-10 z m -2,-12 h 4 l 6,6 h -4 z m -74,28 -4,4 v 10 l 8.12494,8.14285 L 34,296 h 8 v -8 l 6,-6 v -4 l 6,-6 v -4 l 4,-4 v -8 l -4,-4 h -8 l -4,-4 z" clip-path="url(#clipPath987-2)" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.01129821px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:accumulate" transform="matrix(0.96464464,0,0,0.96464464,-475.64889,273.86349)"/>
          <ns0:g transform="matrix(0.33027944,0,0,0.33027944,-722.51179,363.54416)" id="g6008" style="display:inline;opacity:1;stroke:#000000;enable-background:new">
            <ns0:circle r="36.270779" cy="372.21783" cx="883.60425" id="path3066-4" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:16.92636299;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
            <ns0:circle r="68.971695" cy="372.2179" cx="883.60431" id="path3941-2" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:11.69271851;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
            <ns0:circle r="103.1213" cy="372.21796" cx="883.60437" id="path3943-0" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:5.99500418;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
          </ns0:g>
          <ns0:g transform="translate(-477.91161,277.51965)" id="g6092" style="display:inline;enable-background:new">
            <ns0:g id="g6087">
              <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:new" ns2:nodetypes="cccssccc" id="path3970-7-4" d="m 47.589745,209.314 -47.7665216,46.36163 21.7759096,0.70244 c 0,0 -9.131831,18.96611 -9.131831,18.96611 -2.8097966,8.42939 9.834282,11.59041 11.941628,5.26838 0,0 8.42939,-18.96612 8.42939,-18.96612 l 15.453872,16.50755 z" ns1:connector-curvature="0"/>
            </ns0:g>
          </ns0:g>
        </ns0:g>
        <ns0:path style="color:#000000;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:sans-serif;font-variant-ligatures:normal;font-variant-position:normal;font-variant-caps:normal;font-variant-numeric:normal;font-variant-alternates:normal;font-feature-settings:normal;text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;text-decoration-style:solid;text-decoration-color:#000000;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-orientation:mixed;dominant-baseline:auto;baseline-shift:baseline;text-anchor:start;white-space:normal;shape-padding:0;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.7453416;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:new" d="m 618.48523,662.34471 a 1.1180124,1.1180124 0 0 0 -1.11802,1.11801 1.1180124,1.1180124 0 0 0 0.74535,1.05269 v 6.09339 a 1.1180124,1.1180124 0 0 0 -0.74535,1.05268 1.1180124,1.1180124 0 0 0 1.11802,1.11802 1.1180124,1.1180124 0 0 0 0.96716,-0.55901 h 6.26498 a 1.1180124,1.1180124 0 0 0 0.96661,0.55901 1.1180124,1.1180124 0 0 0 1.11802,-1.11802 1.1180124,1.1180124 0 0 0 -0.74535,-1.05268 v -6.09339 a 1.1180124,1.1180124 0 0 0 0.74535,-1.05269 1.1180124,1.1180124 0 0 0 -1.11802,-1.11801 1.1180124,1.1180124 0 0 0 -1.10109,0.93168 h -5.99548 a 1.1180124,1.1180124 0 0 0 -1.10218,-0.93168 z m 0.96716,1.67702 h 6.26498 a 1.1180124,1.1180124 0 0 0 0.0244,0.0426 l -0.96607,0.96607 a 0.74534162,0.74534162 0 0 0 -0.32772,-0.077 0.74534162,0.74534162 0 0 0 -0.7206,0.559 h -2.28497 a 0.74534162,0.74534162 0 0 0 -0.72114,-0.559 0.74534162,0.74534162 0 0 0 -0.32809,0.0766 l -0.96643,-0.96644 a 1.1180124,1.1180124 0 0 0 0.0257,-0.0419 z m -0.59449,0.52698 1.11946,1.11947 a 0.74534162,0.74534162 0 0 0 -9.9e-4,0.0306 0.74534162,0.74534162 0 0 0 0.37267,0.64471 v 2.43765 a 0.74534162,0.74534162 0 0 0 -0.37267,0.64435 0.74534162,0.74534162 0 0 0 0.0766,0.32809 l -0.96644,0.96643 a 1.1180124,1.1180124 0 0 0 -0.22819,-0.11118 z m 7.45341,0 v 6.06009 a 1.1180124,1.1180124 0 0 0 -0.22891,0.11045 l -0.96607,-0.96607 a 0.74534162,0.74534162 0 0 0 0.077,-0.32772 0.74534162,0.74534162 0 0 0 -0.37267,-0.64472 v -2.43764 a 0.74534162,0.74534162 0 0 0 0.37267,-0.64435 0.74534162,0.74534162 0 0 0 -10e-4,-0.0309 z m -5.09838,1.70905 h 2.74299 a 0.74534162,0.74534162 0 0 0 0.11937,0.0857 v 2.43765 a 0.74534162,0.74534162 0 0 0 -0.34793,0.45801 h -2.28497 a 0.74534162,0.74534162 0 0 0 -0.34847,-0.45838 v -2.43764 a 0.74534162,0.74534162 0 0 0 0.11901,-0.0853 z m 0,3.7267 h 2.74299 a 0.74534162,0.74534162 0 0 0 0.49204,0.18634 0.74534162,0.74534162 0 0 0 0.0309,-10e-4 l 1.14349,1.14349 a 1.1180124,1.1180124 0 0 0 -0.0395,0.16195 h -5.99548 a 1.1180124,1.1180124 0 0 0 -0.0411,-0.16141 l 1.1444,-1.14439 a 0.74534162,0.74534162 0 0 0 0.0306,10e-4 0.74534162,0.74534162 0 0 0 0.49168,-0.18634 z" id="path1558" ns1:connector-curvature="0"/>
        <ns0:g transform="matrix(0.0931677,0,0,0.0931677,616.58763,660.31823)" style="display:inline;enable-background:new" id="g1207">
          <ns0:rect ry="8.555583" rx="8.555583" y="176.2498" x="16.944288" height="115.50041" width="94.111382" id="rect15435-6" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:4;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
          <ns0:path style="display:inline;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.0119126px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" d="m 525,430.125 c -2.216,0 -4,1.784 -4,4 V 463 h 80 v -28.875 c 0,-2.216 -1.784,-4 -4,-4 z M 521,465 v 30 h 80 v -30 z m 0,32 v 29 c 0,2.216 1.784,4 4,4 h 72 c 2.216,0 4,-1.784 4,-4 v -29 z" transform="translate(-497,-247)" id="rect15441-8" ns1:connector-curvature="0" ns2:nodetypes="ssccsssccccccsssscc"/>
          <ns0:g id="g1088">
            <ns0:path style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.01184966px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" d="m 552,443 c -1.662,0 -3,1.338 -3,3 v 4 1 h 4 0.0312 l -0.0156,-2 H 569 v 2 H 569.0312 573 v -1 -4 c 0,-2 -1.338,-3 -3,-3 z" transform="translate(-497,-247)" id="path26035" ns1:connector-curvature="0"/>
          </ns0:g>
          <ns0:use height="100%" width="100%" transform="translate(0,32)" id="use1090" ns4:href="#g1088" y="0" x="0"/>
          <ns0:use x="0" y="0" ns4:href="#g1088" id="use1092" transform="translate(0,64)" width="100%" height="100%"/>
        </ns0:g>
        <ns0:g style="display:inline" transform="matrix(0.0931677,0,0,0.0931677,544.00999,756.23256)" id="g16105">
          <ns0:path ns1:connector-curvature="0" id="rect854" d="m 798.33622,-694.6285 c -4.70031,0 -8.48432,3.78401 -8.48432,8.48432 v 10.60536 74.23787 8.48433 c 0,4.70031 3.78401,8.48432 8.48432,8.48432 h 93.32756 c 4.70031,0 8.48432,-3.78401 8.48432,-8.48432 v -8.48433 -74.23787 -10.60536 c 0,-4.70031 -3.78401,-8.48432 -8.48432,-8.48432 z" style="display:inline;opacity:1;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:4;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
          <ns0:rect style="display:inline;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.01121096px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" id="rect858" width="96" height="87.999969" x="797" y="599.48041" rx="4" ry="3.9999695" transform="scale(1,-1)"/>
          <ns0:g style="display:inline;fill:#ffffff;enable-background:new" transform="translate(779,-877.48042)" id="g866">
            <ns0:path ns1:connector-curvature="0" id="path862" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:medium;line-height:1.25;font-family:'Source Code Pro';-inkscape-font-specification:'Source Code Pro, Bold';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.24999999" d="M 44.012301,210.88755 30,203.27182 V 208 l 9.710724,4.62951 v 0.1422 L 30,218 v 4.72818 l 14.012301,-8.21451 z" ns2:nodetypes="ccccccccc"/>
            <ns0:path ns2:nodetypes="ccccc" ns1:connector-curvature="0" id="path864" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:medium;line-height:1.25;font-family:'Source Code Pro';-inkscape-font-specification:'Source Code Pro, Bold';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.24999999" d="m 47.999998,226 2e-6,4 h 16.00001 l -2e-6,-4 z"/>
          </ns0:g>
        </ns0:g>
      </ns0:g>
      <ns0:g id="g1220" style="display:inline" transform="matrix(1.0281734,0,0,1.0281734,706.43823,751.89837)" ns1:label="#g5607">
        <ns0:path d="M 27.135224,2.8483222 V 19.288556 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path1214" style="color:#000000;display:block;overflow:visible;visibility:visible;opacity:0.6;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;filter:url(#filter5601);enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path1216" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient5176);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path d="M 26.604893,2.3179921 V 18.758225 l 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 h 4.684582 z" id="path1218" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient5885);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:rect y="700.19403" x="521.92926" height="3.3540373" width="29.813665" id="rect5339" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle r="4.2555118" cy="701.69794" cx="511.71103" id="circle5343" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.37267077;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect5345" width="28.03303" height="3.3540373" x="521.92926" y="715.10089"/>
      <ns0:rect y="715.10089" x="552.86096" height="3.3540373" width="20.124224" id="rect5347" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5349" cx="511.71103" cy="716.6048" r="4.2555118"/>
      <ns0:rect y="730.00775" x="521.92926" height="3.3540373" width="25.341616" id="rect5351" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle r="4.2555118" cy="731.51166" cx="511.71103" id="circle5355" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect5357" width="17.888199" height="3.3540373" x="521.92926" y="744.91461"/>
      <ns0:rect y="744.91461" x="544.28955" height="3.3540373" width="28.695652" id="rect5359" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle5361" cx="511.71103" cy="746.41852" r="4.2555118"/>
      <ns0:rect y="759.82147" x="521.92926" height="3.3540373" width="30.931677" id="rect5363" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle r="4.2555118" cy="761.32538" cx="511.71103" id="circle5367" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:g style="display:inline;stroke:#ffffff;enable-background:new" id="g2204" ns1:label="edit-find" transform="matrix(0.37267081,0,0,0.37267081,456.52122,410.84515)">
        <ns0:circle transform="matrix(1.2871768,0,0,1.2857143,-249.29926,155.57143)" id="path27918" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#ffffff;stroke-width:1.55467153;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" cx="307.5" cy="386.5" r="3.5"/>
        <ns0:path ns2:nodetypes="cc" id="path27941" d="m 150.01159,656.00001 4.00455,4" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#ffffff;stroke-width:2;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" ns1:connector-curvature="0"/>
      </ns0:g>
    </ns0:g>
  </ns0:g>
</ns0:svg>
