<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Byt skrivbordsbakgrund</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="prefs-display.html" title="Visning och skärm">Visning och skärm</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Byt skrivbordsbakgrund</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan ändra vilken bild som används som skrivbordsbakgrund, eller använda en enkel färg eller färgskala.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Högerklicka på skrivbordet och välj <span class="gui">Byt skrivbordsbakgrund</span>.</p></li>
<li class="steps"><p class="p">Select an image or color. The settings are applied immediately.
  <span class="link"><a href="shell-workspaces-switch.html" title="Switch between workspaces">Switch to an empty workspace</a></span>
  to view your entire desktop.</p></li>
</ol></div></div></div>
<p class="p">Det finns tre val i den utfällbara listan längst upp till höger.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list">
<p class="p">Välj <span class="gui">Bakgrundsbilder</span> för att använda en av de många bilder som skapats av yrkeskunniga som distribueras tillsammans med Ubuntu. Med undantag för Ubuntus bakgrundsbild skapades alla standardbakgrunder av vinnarna av en skrivbordsbakgrundstävling inom gemenskapen.</p>
<p class="p">Vissa bakgrundsbilder är delvis genomskinliga och tillåter att en bakgrundsfärg syns igenom. För dessa skrivbordsbakgrunder kommer det finnas en färgvalsknapp längst ner till höger.</p>
</li>
<li class="list"><p class="p">Välj <span class="gui">Bildmapp</span> för att använda en av dina egna bilder från din Bildmapp. De flesta bildhanteringsprogram lagrar foton där.</p></li>
<li class="list"><p class="p">Välj <span class="gui">Färger &amp; tonskalor</span> för att bara använda en enkel färg eller en linjär färgtonskala. Färgvalsknappar kommer visas längst ner till höger.</p></li>
</ul></div></div></div>
<p class="p">Du kan också bläddra bland bilderna på din dator genom att klicka på <span class="gui">+</span>-knappen. Bilderna du lägger till på det här sättet kommer visas under mappen <span class="gui">Bilder</span>. Du kan ta bort den från listan genom att markera den och klicka på <span class="gui">-</span>-knappen. Bilder som tas bort från listan kommer inte raderas från disken.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs-display.html" title="Visning och skärm">Visning och skärm</a><span class="desc"> — 
      <span class="link"><a href="look-background.html" title="Byt skrivbordsbakgrund">Background</a></span>,
      <span class="link"><a href="look-resolution.html" title="Ändra storlek och rotation för skärmen">size and rotation</a></span>,
      <span class="link"><a href="display-dimscreen.html" title="Ställ in skärmens ljusstyrka">brightness</a></span>…
    </span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
