<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Tidssynkronisering med NTP</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="networking.html" title="Nätverk">Nätverk</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="dhcp.html" title="Dynamic Host Configuration Protocol (DHCP)">Föregående</a><a class="nextlinks-next" href="DPDK.html" title="Data Plane Development Kit">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Tidssynkronisering med NTP</h1></div>
<div class="region">
<div class="contents">
<p class="para">NTP är ett TCP/IP protokoll för synkronisering av tid över ett nätverk. I grund och botten är det en klient som frågar en server efter nuvarande tid och använder det för att ställa in sin egen klocka.</p>
<p class="para">
Behind this simple description, there is a lot of complexity - there are tiers of NTP servers, with the tier one NTP servers connected to atomic clocks, and tier two and three servers spreading the load of actually handling requests across the Internet. Also the client software is a lot more complex than you might think - it has to factor out communication delays, and adjust the time in a way that does not upset all the other processes that run on the server. But luckily all that complexity is hidden from you! 
</p>
<p class="para">
Ubuntu uses ntpdate and ntpd. 
</p>
</div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="NTP.html#timedatectl" title="timedatectl">timedatectl</a></li>
<li class="links"><a class="xref" href="NTP.html#timesyncd" title="timesyncd">timesyncd</a></li>
<li class="links"><a class="xref" href="NTP.html#ntpdate" title="ntpdate">ntpdate</a></li>
<li class="links"><a class="xref" href="NTP.html#timeservers" title="timeservers">timeservers</a></li>
<li class="links"><a class="xref" href="NTP.html#ntpd" title="ntpd">ntpd</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-installation" title="Installation">Installation</a></li>
<li class="links"><a class="xref" href="NTP.html#timeservers-conf" title="Konfiguration">Konfiguration</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-status" title="View status">View status</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-pps" title="PPS Support">PPS Support</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-references" title="Referenser">Referenser</a></li>
</ul></div>
<div class="sect2 sect" id="timedatectl"><div class="inner">
<div class="hgroup"><h2 class="title">timedatectl</h2></div>
<div class="region"><div class="contents">
<p class="para">
		In recent Ubuntu releases <span class="em emphasis">timedatectl</span> replaces <span class="em emphasis">ntpdate</span>.
		By default <span class="em emphasis">timedatectl</span> syncs the time once on boot and later on uses socket activation to recheck once network connections become active.
</p>
<p class="para">
		If <span class="em emphasis">ntpdate / ntp</span> is installed <span class="em emphasis">timedatectl</span> steps back to let you keep your old setup.
		That shall ensure that no two time syncing services are fighting and also to retain any kind of old behaviour/config that you had through an upgrade.
		But it also implies that on an upgrade from a former release ntp/ntpdate might still be installed and therefore renders the new systemd based services disabled.
</p>
</div></div>
</div></div>
<div class="sect2 sect" id="timesyncd"><div class="inner">
<div class="hgroup"><h2 class="title">timesyncd</h2></div>
<div class="region"><div class="contents">
<p class="para">
		In recent Ubuntu releases <span class="em emphasis">timesyncd</span> replaces the client portion of <span class="em emphasis">ntpd</span>.
		By default <span class="em emphasis">timesyncd</span> regularly checks and keeps the time in sync.
		It also stores time updates locally, so that after reboots monotonically advances if applicable.
</p>
<p class="para">
		The current status of time and time configuration via <span class="em emphasis">timedatectl</span> and <span class="em emphasis">timesyncd</span> can be checked with <span class="em emphasis">timedatectl status</span>.
</p>
<div class="code"><pre class="contents ">timedatectl status
      Local time: Fri 2016-04-29 06:32:57 UTC
  Universal time: Fri 2016-04-29 06:32:57 UTC
        RTC time: Fri 2016-04-29 07:44:02
       Time zone: Etc/UTC (UTC, +0000)
 Network time on: yes
NTP synchronized: no
 RTC in local TZ: no
</pre></div>
<p class="para">
		If NTP is installed and replaces the activity of <span class="em emphasis">timedatectl</span> the line "NTP synchronized" is set to yes.
</p>
<p class="para">
		The nameserver to fetch time for <span class="em emphasis">timedatectl</span> and <span class="em emphasis">timesyncd</span> from can be specified in /etc/systemd/timesyncd.conf and with flexible additional config files in /etc/systemd/timesyncd.conf.d/.
</p>
</div></div>
</div></div>
<div class="sect2 sect" id="ntpdate"><div class="inner">
<div class="hgroup"><h2 class="title">ntpdate</h2></div>
<div class="region"><div class="contents">
<p class="para">
		<span class="em emphasis">ntpdate</span> is considered deprecated in favour of <span class="em emphasis">timedatectl</span> and thereby no more installed by default.
		If installed it will run once at boot time to set up your time according to Ubuntu's NTP server.
		Later on anytime a new interface comes up it retries to update the time - while doing so it will try to slowly drift time as long as the delta it has to cover isn't too big.
		That behaviour can be controlled with the <span class="em emphasis">-B/-b</span> switches.
</p>
<div class="code"><pre class="contents ">ntpdate ntp.ubuntu.com
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="timeservers"><div class="inner">
<div class="hgroup"><h2 class="title">timeservers</h2></div>
<div class="region"><div class="contents"><p class="para">
	   By default the systemd based tools request time information at ntp.ubuntu.com.
	   In classic ntpd based service uses the pool of [0-3].ubuntu.pool.ntp.org
	   Of the pool number 2.ubuntu.pool.ntp.org as well as ntp.ubuntu.com also support ipv6 if needed.
	   If one needs to force ipv6 there also is ipv6.ntp.ubuntu.com which is not configured by default.
   </p></div></div>
</div></div>
<div class="sect2 sect" id="ntpd"><div class="inner">
<div class="hgroup"><h2 class="title">ntpd</h2></div>
<div class="region"><div class="contents"><p class="para">
   The ntp daemon ntpd calculates the drift of your system clock and continuously adjusts it, so there are no large corrections that could 
   lead to inconsistent logs for instance. The cost is a little processing power and memory, but for a modern server this is negligible. 
   </p></div></div>
</div></div>
<div class="sect2 sect" id="ntp-installation"><div class="inner">
<div class="hgroup"><h2 class="title">Installation</h2></div>
<div class="region"><div class="contents">
<p class="para">
   To install ntpd, from a terminal prompt enter: 
   </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install ntp</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="timeservers-conf"><div class="inner">
<div class="hgroup"><h2 class="title">Konfiguration</h2></div>
<div class="region"><div class="contents">
<p class="para">
  Edit <span class="file filename">/etc/ntp.conf</span> to add/remove server lines.
  By default these servers are configured:
  </p>
<div class="code"><pre class="contents "># Use servers from the NTP Pool Project. Approved by Ubuntu Technical Board
# on 2011-02-08 (LP: #104525). See http://www.pool.ntp.org/join.html for
# more information.
server 0.ubuntu.pool.ntp.org
server 1.ubuntu.pool.ntp.org
server 2.ubuntu.pool.ntp.org
server 3.ubuntu.pool.ntp.org
</pre></div>
<p class="para">
	  After changing the config file you have to reload the
          <span class="app application">ntpd</span>:
	  </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo systemctl reload ntp.service</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="ntp-status"><div class="inner">
<div class="hgroup"><h2 class="title">View status</h2></div>
<div class="region"><div class="contents">
<p class="para">
  Use ntpq to see more info: 
  </p>
<div class="screen"><pre class="contents "><span class="cmd command"># sudo ntpq -p</span>
<span class="output computeroutput">     remote           refid      st t when poll reach   delay   offset  jitter
==============================================================================
+stratum2-2.NTP. 129.70.130.70    2 u    5   64  377   68.461  -44.274 110.334
+ntp2.m-online.n 212.18.1.106     2 u    5   64  377   54.629  -27.318  78.882
*145.253.66.170  .DCFa.           1 u   10   64  377   83.607  -30.159  68.343
+stratum2-3.NTP. 129.70.130.70    2 u    5   64  357   68.795  -68.168 104.612
+europium.canoni 193.79.237.14    2 u   63   64  337   81.534  -67.968  92.792</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="ntp-pps"><div class="inner">
<div class="hgroup"><h2 class="title">PPS Support</h2></div>
<div class="region"><div class="contents"><p class="para">
Since 16.04 ntp supports PPS discipline which can be used to augment ntp with local timesources for better accuracy.
For more details on configuration see the external pps ressource listed below.
  </p></div></div>
</div></div>
<div class="sect2 sect" id="ntp-references"><div class="inner">
<div class="hgroup"><h2 class="title">Referenser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
  	    <p class="para">
          See the <a href="https://help.ubuntu.com/community/UbuntuTime" class="ulink" title="https://help.ubuntu.com/community/UbuntuTime">Ubuntu Time</a> wiki page for more information.
        </p>
      </li>
<li class="list itemizedlist">
  	    <p class="para">
          <a href="http://www.ntp.org/" class="ulink" title="http://www.ntp.org/">ntp.org, home of the Network Time Protocol project</a>
        </p>
      </li>
<li class="list itemizedlist">
  	    <p class="para">
		    <a href="http://www.ntp.org/ntpfaq/NTP-s-config-adv.htm#S-CONFIG-ADV-PPS" class="ulink" title="http://www.ntp.org/ntpfaq/NTP-s-config-adv.htm#S-CONFIG-ADV-PPS">ntp.org faq on configuring PPS</a>
        </p>
      </li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="dhcp.html" title="Dynamic Host Configuration Protocol (DHCP)">Föregående</a><a class="nextlinks-next" href="DPDK.html" title="Data Plane Development Kit">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
