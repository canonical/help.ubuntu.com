<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" height="500" id="svg10075" version="1.1" width="840" ns2:docname="gs-goa5.svg" ns1:version="0.92.4 5da689c313, 2019-01-14">
  <ns0:defs id="defs10077">
    <ns0:linearGradient id="RHEL7" ns3:paint="gradient">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop id="stop11074" offset="0" style="stop-color:#eeedec;stop-opacity:1;"/>
      <ns0:stop id="stop11076" offset="1" style="stop-color:#eeedec;stop-opacity:1"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop id="stop7012" offset="0" style="stop-color:#eeedec;stop-opacity:0;"/>
      <ns0:stop id="stop7014" offset="1" style="stop-color:#eeedec;stop-opacity:0"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" gradientUnits="userSpaceOnUse" id="linearGradient7064" x1="-18.33782" x2="713.42853" y1="490.54935" y2="490.54935" ns1:collect="always" ns4:href="#GNOME"/>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient5885" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop id="stop5718" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17441" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop id="stop17445" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop17447" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17453" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17455" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:filter color-interpolation-filters="sRGB" height="1.1308649" id="filter5601" width="1.2058235" x="-0.10291173" y="-0.065432459" ns1:collect="always">
      <ns0:feGaussianBlur id="feGaussianBlur5603" stdDeviation="0.610872" ns1:collect="always"/>
    </ns0:filter>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17453-7" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716-4"/>
    <ns0:linearGradient id="linearGradient5716-4">
      <ns0:stop id="stop5718-1" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720-6" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17455-1" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716-4"/>
    <ns0:linearGradient id="linearGradient16929">
      <ns0:stop id="stop16931" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop16933" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
  </ns0:defs>
  <ns2:namedview bordercolor="#666666" borderlayer="true" borderopacity="1.0" fit-margin-bottom="0" fit-margin-left="0" fit-margin-right="0" fit-margin-top="0" height="0px" id="base" pagecolor="#eeeeec" showgrid="false" width="0px" ns1:current-layer="layer2" ns1:cx="383.02942" ns1:cy="302.54948" ns1:document-units="px" ns1:pageopacity="1" ns1:pageshadow="2" ns1:showpageshadow="false" ns1:window-height="1249" ns1:window-maximized="0" ns1:window-width="1484" ns1:window-x="355" ns1:window-y="132" ns1:zoom="1">
    <ns1:grid empspacing="5" enabled="true" id="grid17504" snapvisiblegridlinesonly="true" type="xygrid" visible="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true" ns1:groupmode="layer" ns1:label="bg">
    <ns0:rect height="656" id="background" style="fill:url(#BLANK);" width="866" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g id="layer2" transform="translate(0,-540)" ns1:groupmode="layer" ns1:label="fg">
    <ns0:g id="g11020" transform="translate(-35,-141.36217)">
      <ns0:circle cx="120" cy="278" id="path11014" r="17" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;enable-background:accumulate" transform="translate(2,453.36217)"/>
      <ns0:text id="text11016" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" xml:space="preserve"><ns0:tspan id="tspan11018" style="font-size:14px;line-height:1.25" x="122.29289" y="736.36218" ns2:role="line">6</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g id="g4890" style="display:inline" transform="matrix(2.6833333,0,0,2.6833333,-1275.5101,-1072.8539)">
      <ns0:g id="default-pointer-c" style="display:inline" transform="matrix(1.0281734,0,0,1.0281734,813.41674,729.17439)" ns1:label="#g5607">
        <ns0:path d="m 27.135224,2.8483222 0,16.4402338 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 27.135224,2.8483222 z" id="path5567" style="opacity:0.6;color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;filter:url(#filter5601);enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path5565" style="color:#000000;fill:url(#linearGradient17453-7);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        <ns0:path d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path6242" style="color:#000000;fill:url(#linearGradient17455-1);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
      </ns0:g>
      <ns0:rect height="168.81989" id="rect4889" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" width="167.70187" x="556.96027" y="608.88965"/>
      <ns0:text id="text26176" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.47858" y="635.46222" xml:space="preserve"><ns0:tspan id="tspan26178" style="font-size:5.21739101px;line-height:1.25" x="610.47858" y="635.46222" ns2:role="line">Google</ns0:tspan></ns0:text>
      <ns0:text id="text26182" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.47858" y="642.17023" xml:space="preserve"><ns0:tspan id="tspan26184" style="font-size:4.47205019px;line-height:1.25" x="610.47858" y="642.17023" ns2:role="line">maria.johansson@gmail.com</ns0:tspan></ns0:text>
      <ns0:text id="text26186" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="611.59662" y="666.76648" xml:space="preserve"><ns0:tspan id="tspan26188" style="font-size:5.21739101px;line-height:1.25" x="611.59662" y="666.76648" ns2:role="line">Använd för</ns0:tspan></ns0:text>
      <ns0:text id="text26190" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="666.76648" xml:space="preserve"><ns0:tspan id="tspan26192" style="font-size:5.21739101px;line-height:1.25" x="622.40393" y="666.76648" ns2:role="line">E-post</ns0:tspan></ns0:text>
      <ns0:text id="text28655" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="679.43726" xml:space="preserve"><ns0:tspan id="tspan28657" style="font-size:5.21739101px;line-height:1.25" x="622.40393" y="679.43726" ns2:role="line">Kalender</ns0:tspan></ns0:text>
      <ns0:text id="text28673" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="692.10803" xml:space="preserve"><ns0:tspan id="tspan28675" style="font-size:5.21739101px;line-height:1.25" x="622.40393" y="692.10803" ns2:role="line">Kontakter</ns0:tspan></ns0:text>
      <ns0:text id="text28691" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="704.77881" xml:space="preserve"><ns0:tspan id="tspan28693" style="font-size:5.21739101px;line-height:1.25" x="622.40393" y="704.77881" ns2:role="line">Foto</ns0:tspan></ns0:text>
      <ns0:text id="text28709" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="717.44958" xml:space="preserve"><ns0:tspan id="tspan28711" style="font-size:5.21739101px;line-height:1.25" x="622.40393" y="717.44958" ns2:role="line">Filer</ns0:tspan></ns0:text>
      <ns0:rect height="10.92049" id="rect3923-9" rx="5.4602423" ry="5.4602423" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" width="19.803892" x="670.62494" y="660.20514"/>
      <ns0:circle cx="684.57684" cy="665.66193" id="path915" r="4.4139271" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:path d="m 600.84504,636.65363 a 5.3133016,5.3133016 0 0 1 -3.93812,5.13225 5.3133016,5.3133016 0 0 1 -5.97664,-2.4756 5.3133016,5.3133016 0 0 1 0.84439,-6.41373 5.3133016,5.3133016 0 0 1 6.41372,-0.84438" id="path4883" style="opacity:1;vector-effect:none;fill:none;fill-opacity:1;stroke:#000000;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" ns2:cx="595.53174" ns2:cy="636.65363" ns2:end="5.2359878" ns2:open="true" ns2:rx="5.3133016" ns2:ry="5.3133016" ns2:start="0" ns2:type="arc"/>
      <ns0:path d="m 595.9382,635.63421 v 2.53516 h 5.48321 l 0.69267,-1.30041 0.0155,-1.23475 z" id="path4885" style="color:#000000;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:sans-serif;font-variant-ligatures:normal;font-variant-position:normal;font-variant-caps:normal;font-variant-numeric:normal;font-variant-alternates:normal;font-feature-settings:normal;text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;text-decoration-style:solid;text-decoration-color:#000000;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-orientation:mixed;dominant-baseline:auto;baseline-shift:baseline;text-anchor:start;white-space:normal;shape-padding:0;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" ns2:nodetypes="cccccc" ns1:connector-curvature="0"/>
      <ns0:rect height="10.92049" id="rect4891" rx="5.4602423" ry="5.4602423" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" width="19.803892" x="670.62494" y="672.8761"/>
      <ns0:circle cx="684.57684" cy="678.33289" id="circle4893" r="4.4139271" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect height="10.92049" id="rect4899" rx="5.4602423" ry="5.4602423" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" width="19.803892" x="670.62494" y="685.54669"/>
      <ns0:circle cx="684.57684" cy="691.00348" id="circle4901" r="4.4139271" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect height="10.92049" id="rect4903" rx="5.4602423" ry="5.4602423" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" width="19.803892" x="670.62494" y="698.21765"/>
      <ns0:circle cx="684.57684" cy="703.67444" id="circle4905" r="4.4139271" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect height="10.92049" id="rect4907" rx="5.4602423" ry="5.4602423" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" width="19.803892" x="670.62494" y="710.88824"/>
      <ns0:circle cx="684.57684" cy="716.34503" id="circle4909" r="4.4139271" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect height="10.92049" id="rect4911" rx="5.4602423" ry="5.4602423" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708" width="19.803892" x="670.62494" y="723.5592"/>
      <ns0:circle cx="684.57684" cy="729.01599" id="circle4913" r="4.4139271" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:text id="text4917" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="622.40393" y="730.86591" xml:space="preserve"><ns0:tspan id="tspan4915" style="font-size:5.21739101px;line-height:1.25" x="622.40393" y="730.86591" ns2:role="line">Skriv­ar­e</ns0:tspan></ns0:text>
      <ns0:rect height="16.397507" id="rect4919" rx="2.9813664" ry="2.9813664" style="opacity:1;vector-effect:none;fill:#c01c28;fill-opacity:1;stroke:none;stroke-width:2.53416157;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" width="54.782524" x="659.81744" y="750.8772"/>
      <ns0:text id="text4923" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.46583843px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.3726708" x="666.71997" y="760.92218" xml:space="preserve"><ns0:tspan id="tspan4921" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.46583843px;font-family:Cantarell;-inkscape-font-specification:Cantarell;fill:#ffffff;stroke-width:0.3726708" x="666.71997" y="760.92218" ns2:role="line">Ta bort konto</ns0:tspan></ns0:text>
    </ns0:g>
  </ns0:g>
</ns0:svg>
