�PNG

   IHDR  !  �   W5"w   �zTXtRaw profile type exif  x�mP[!��=�<t�8n�&�A�_Lv۝�a�8"�?�<$o�h)� *J�DM�6�L� ��:��,�e�F-�q�����L��3�����x��Dd�##&o`4�V*Z������0h�9Q�?�f�;���D���Y| ���ہ��8Ge��r����jZ�3fL  �iCCPICC profile  x�}�=H�@�_S�"�q�P����U(B�P+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�F�iV�,�鶙N&�lnU�"�D0Qf�1'I)���{�z�Y���}j�b@@$�e�ioOo��}�(+�*�9�I$~�����ό���<q�X,v����dj�S�1U�)_�z�r��Uj�uO��p^_Y�:�a$��%H���2*��U'�B��>�!�/�K!W��B������w�Var�K
'����B�@��8�ǎ�<������W��'���;����붦��;���!��+i
��~Fߔ"�@��[k�@��J� ��h���}����ۿgZ�� ��r�(˞�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:366edc7c-fd23-4cb7-875c-39ca03d3db38"
   xmpMM:InstanceID="xmp.iid:cf7c2a01-7117-482f-b9ec-3771b8fc2d58"
   xmpMM:OriginalDocumentID="xmp.did:5060ddc3-8834-4dbf-be28-4544e7b41613"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679601200580845"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T20:53:20+01:00"
   xmp:ModifyDate="2023:03:23T20:53:20+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:7191b091-720c-4ac1-a830-13d0a22d6403"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T20:53:20+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>�Ѕ   	pHYs  �  ��+   tIME�
*==   tEXtComment Created with GIMPW�    IDATx��wt\�u.���w� 0轱��"Ţ�H[5�mI.�Ǳ���V���;���ʎc'�$ۊ%Q�*I�EI��" ���`�ܳ�{	� g@����-��;�ܲ����go��@BbP�����t�JD�)HHL�|R�Iܒ���s䃐�4��g  �|�E�	�%��f���c'["}>��秫��[-& �s]����s_�v�������?<�K���Ĕ�Lex�,��9ݪIA_��wD������D�>'���w� P}1|M[Tb�8k��*��_�
:-,;U���Ӿ�BW���!�\�6� �HpΛ��/^��06}����L �p�bsS��yyYYaa!c�DQKK�� `ZUUvv6"�b��������¢��EQ.�֐�_{��ܹs�V+缶����3;;{��pyW�y�濹Ǖbe�y��-)����i���w"�LU@1��b?��,��~8�?���T3r�Qm[t�o��J/r�?�9�`V����}���΁�q����D�������?��/j��9�����A_ww����mkkkrG�B�7����W[[��/":~���m�����������֛o���+|>UWW���n x��9rc_M��mK��p�~�k��6{w�	@U�i^�y"T
Q��!���	V�V�u�+;U�������e(�=N�a��&?�<�*���~�P\}~�҇C�K,�.p��*zLڊ7��i_�����������p8l��>��? M�/��7��䋃[ZZ��p__��f���mkkG�e��iii=^osSs,+**����4���<2�BU�U˰�ڬ�o|��88����/>ߠɤ����>�LQaQV�g��Θ1}�k[E���uDT}�f�7���$�P(���w���gsrrfΘ�a�ƙ3����$%�Q�m����G� ��Ђ"K���Mȼ�S\����������_�������`Z���Ģ�*�p`(�����L��g�s���|o���3y0J�k��vv�l�����Ψ��n�x������_Ӵ��������޽{�[[�*+O�:m�Z����Z[�����p���������;w�������s�UTTTUU����ͦ+G�F#��*�������� �������9�;w"���رcw�\��׀H�b�X�����9�Ή��W�� �L������k��&��ڰv�:5ө���<8�>;xZ��ߨ��|si�ǞL�v�%�����{cDֱΜT%����@so��l��� `���ӟJq;����n.��СCӧM3�T �ny�����f��̤ys��s�]EE�;w�����wvv��׿��ϟW\\�������[Z����n��u��/�9������ljn6�L�0���F����\P��]��O�VXX��A�m�ܹ�lذxѢ�3gb1-�&�9l?XTb�LQ~�yO��Wd�f��'[��|+ϥ�-�d�*�Z# p�9 �n57Mq�ؙ��E�*p�8A��x�G��D4L���N��hQ�o2�m8w���/|�Y�:l6�g������mݺuǎ��>�t<d�**"z2=�5;���ڡ�G�.5���9�h$JD��Z,q�+Gljj޿��3O�d29��@0�FUUC6���ↆso��μ�sO~��ٳg���K_���{>�����ٳg����͖���Վ��\�����˭٩�p�4��zƋ+���}�[�|�S)����Ե�m�}����m����JV�2;�|�)l5����y��>�7���X�>���RK�O��k��c�b7�Jl8װa�?y����"��mV��l���=w�q��P�࢑�W ػw�c�<RXXx�S@@@4�X��_��{����┙��JM=~��ܹs
��7�B�իW�����(
utt�Y��j�Fc�eK��'R�����	��U�8��3貱9�f �����ۧ��H[5�洲�����;��{q��n��<���7�Fe���_��S�e��թ��& `-}�׎�Ť`�������ы��/wz��G-��F[]�8��荍��$�n }������v������e˲��6m�L�Y�=w�#��� �@��l...ڲu[^^���k&����H$��_�'~��ѣ55�6s�����w�9y�ohh��#bII	2�٬��< �v�=77>|����d6�B���̦֙	�]�������ֻ�2��O�Q�q#��t;�Yy��n�`	 ��7�l�[�1N��Z����q@So�o7���}_���?L��w�;�v��u���iy.ei��L{��C��x׌}=]R�o��hùsd,v��祦�vww� @zZzFf�b8T===&���r�#������\�im��~����]UT���v��K[[{Vv��d�����?˹.=�9ٙ睝�C�!w�;���+�	�y{{GVv����}}]��
c���rM�f�t�7^���KJ,���>���?�e�?|%K���l�6 o}3GB8�W�-��1Gxh��?��5���L�qǮB�tu�t�3�N�9��[�}&x�e�����on�&���-rL�1�?�7�����S�2T ���ˇ�&�\v��ݝR$&�c]��-1�T�ILV�G>�1�Ab�H&EK�1� $$�&�ր��'Y�������#�A`|B#?��K"�Da����ď�g��J��				>~_�wL֫G�Z��.���3>	��e�B{ W��cG}����+�<�)��.��UD�c;<���~�8��j�W����u�M���	0'�V�(��*ϓ.��Q���2��C@��!�H��q$D" B $�MD�����HH@�8p �\�@ ��� p���/�P?!#�eH#��#!!C�2�=�иr1��7�@�Hd�]� �� �8 
��"�s� G�z�P8p}/��@"@"�o��Ⳍ���4,�\g:h@�#�4�e�hq:���x>��h����I�\����t<q�	9!ň��#�X�f� ��h�/��������"�& D��@4�@ Q�R�0D���E�?{�f�����t�6 ҟ'��c��G|qļG�s�H@@�鯛 8E	��8�s����l ND������	T1�!1]<Q�#��Ef$�߳X�qd@b�� I�'@�!pqR�%_�'�sЙ�s�ǥ�!S�H|�"�t-�8p@f\3
�&�U�rC�q1��:�����@#��3V!��-���0}��/���ڸ� C{�O���>	2s�'1�ǒNeD}b L�[Ɖ��(4��7�c��4��ĭ&0`b�8뙸I4�q1@��[�� '���FX#�W�<�OY�m�%$P'���3��3}�ŏӏИ�I�� F �� ��1��54���� ���pZ�Β�u��g�� �0щ�<7,fj��p�Ft���  r�@#��CRp�0CǠ��9h�Ā�
#Q����j8Gȁ����p5Q���3��I��H���7"��}@ �s���^H@�8Gd��%�`��j�
B�� ���Y�����X�H�D���Jq��P׮\��uA%)� �,�8qa���(&1����^�af�W7"��t(Θ�Wn@";]Lm�z���N������3��i�>1�# B`@�?3�fh���)�9��fc@�17na������_�P_#�"��D�2"�	�#�L�v�O,\(���Awi@L�����G�}D�G"�'�]��Z$b�:1EQ�R-�����y���gD��\���M#'��r ML�q�S(4�D������>ˁ ��xB�\<eÌ��"�3�,��u�
�۲����x�����Y�tfq4�jD ��K- �8�f��%!��i�9#D��A���1(��i�^�0Eㆪn2��IW��nC�	Z|�Ѹ�aJb����[t��y'�1}���ō���qO
8
2"l����
�9�t3[�a �kB`��%�C�[h�Hd���
�AL�������x*�@cz����)q $�8R��W�S���U30E8P7C�R�.���(�����@W���m��������dD􉖄�a`�qr8�$Ll@U�@B�0�@��i� T�� 1e��1E��B�0��v`��"��\�8�[+�X��n[iy�|�n��������q������y6���F�X5 >��?��i7����8aPI��F@'��eӘ�1 ���c\K����:��}��} �	kY'�sø����`@eN��"�4L?aHc���� q�)Ī�,�U� ����zCPU���:}f��e���8���:\�t� ��*^���u���?1Vb�qnvh3�����b��K��Y��wWT���^��	�HV|ˈ��1|D ev�:�L �^,���#lK��@s���,=�IOK���Nk��<�Imm�F5-ݏ/��u�2��a# �#$����rwN_��)$�H|¡(��(�ᰵ��F"���$Ȍe2ev����B����b��XQ-�|� �fdd:�uD�1F#4��|L��G"$}��� �g�bK���)�Iڇ� ��g䯹s��b6�1�"��@P�<���#�3v@d�q���Ӝ����e�CB�J���0SQ�\C���"V�X<��	\��#�"+�8qn�R��d����g�t�����#E�1�b�1�`�F�/h�,#$�$$Ɓ٤���m��N������Hg�]-F��4���W^�I)!!q�c����`Q��Fd9�R��%1}_Jq�
/�����U����r���+B����7|,��!}��c 2�Zㆩ�1X�|z���wH�z��L�]�0 c�"���S2�d��T~��Ή8���n�(-M�)�	>�9��d�s��h�F�G2,��t,�Y�8�kh�o��e/���K
x
���un�4�5>~�+�H�kqJd�acIL����5�j�QpC�	l�챈�����5"� 8#$��l��9S!��œ�'6=p-�M��h��5~�n�X�H0N��9���ȵk{�7x�t���2ox�'R|����2\�%5-�kz�s�z&a�]�Wn�X�J0ε�����Krǚ�M&��4�l6��f����D(��iYE
MX9�DdW��7�X�j"j�23�i��6�v-c��f[m&1��91B�#��n�T�.�h�^�#���\cIL�K�n'�	
Í \i��t�p�D �Qh��8�Łf�D��xDVؾ7�X��d���9��@�+�^pP�~�FP�X�j����7䫫;
��f͜���>�D����%]�]��gK���v��%1�*��% N�`�c�9s&555///��F��q�� TALq#�Z�b�O��lM��~ 8R]���f6���hkk��e�\.���PUuT+Ǯ5�,:;:S]�555��u��-))N��`FFfJJ�X#�JUSD��B8>]{�̙z��<w�܊��q֩��8U��+����:�#�G�J��v;�R]���k�� $�A��.^� ^� �+=F1�q�5����۱s�ѣG5��]�v��5���������g�@NN�hw�8����cEc�~�o߾�����N ��|uuuug��������ƒ�dOl|��;V]}4/77��Nמ���k��_$�=�3V$=q�Įݻ��Қ����Қ[Z�>��Ju���c��c ���C�hlwV	GS' B��t�2!���TW����w�}�p�⥣Gk���V�Z����s5ǎ͜9��p�v�k�!c�q�y���n����?����9EU�>�Ĕ豫�u���+W���۶m=��0���v�Ʊ.]�X}�z��ye���} �.��߳go~^��j�ֱF���l2*������s��-bv�	�cc�a���ܜ��̓'N֝�s8�m��:�t:�����!�k�^�8�?�X}}}��P^^��c�?p�O<��ܹscCC~o�wt(��L����P0%5�l6����L�p(tU�^�XǏ�x<�-�X,6��l6���}�������:�	UU��tTD��pY��<�!����+W��1cFGg�-[���M�[n�s�����ع����d2UVT��v PuZմ��Ʈ����y��'��'>�Ĥ"���d$���mkk ��������O��6��s����Z�t��#֬Y#W���r�vuu%>�HCPn�\4׹�WB�čäH�8�Lv���䢣�������������C��Ν;�*���<#{�YYY�� D����1�Q�&Q�4y�N�����ȑ#�lg׮]�9����ⵎr�=w���F�цs�@  4M������O����7�m-���M�4m'B~J�� @vvNKKK,�aoo���`vvV�c��G ��F݀b�&|�����!�b��l^�f�ɏ>jnn.*,Z�xQ�3����16������+==ݕ����F�כ���������9w:�C���U%�*3(�) x=c�6��ww:th޼yv��s������q挙�c5].\��ո����ĉ��է5˓U�~�?Đ�'3 �����.�;c�x�8��8c��@�PUվ�>ac�LfD��4M3�&��n"����ǆg����ŋ>|���%33SӴ��v\�j��b���F1�ߧ�7�9���g<	C�F9|ժ;���t�ҕ�gZZ��U�G��p���c�e2��.]Z\\�Js>t���6?/�����ȴZ�c�j�fS��p,�9��ܼP��@�8�c��q�2�L�����d�9s���KQԊ��ٳg���^�X��d�EK_�+DD�H#�)�_�����eD�ŒV�TQ��s��:VWWWCCCAAA�TWKbA�iZ��~�S�M1�x��|��n@E  N��tV""ä���S%8VVVV<F��X�j,�e�\���U���2��Fz�zG$4ҩ�M��$���q#ǒ�<0���	�F��]Un�XWGt�1�r��,ѵNK,�>���cIL�W��[@�	��F��q���0BDF��f����9��$rQQ�uK>2T&�o�X#�ӌm���Į]v����u��9�ĤҌ)�u���Z�,�8�m!�^� T F����uxeql��L��__��F�%1��L�	�hA�މ�F� �` T�ȍ�uz���~d��9���%X��F�%1�4CET��q��bm
�o�X�E$TE7[BNH�!�#���j�K�d��o�X��.��Z��M���X�M P	�"�gQ�-k�0?�(�!w4���?��@C��:gz�?�Q%_��D��h��UQ��G ג,!!q���pZH}4u���Hf���H�f�(���H�����DB# ���
3���^��H�C���_� ��IRc���D\l%� z?h�OB"1а2�  0[�YR���6���refd���Z�V���U,���	��H8������	C�p8�m�FmB U/F��w��KV	EQrsr�rssr��6�|�7?<�L �i��������!�?�S���H*  !�D�bJ(,��VU���c��囓���*�Ǔ�v����ן=��|yq�k#��*jx��N\���1�I-*(�7w��,�%qCQWj�r��O��^����ĉ!�(2@H9��T�V���RL����Ens��^����@����E D��r���Ι5sάY�`L@�,�g���n�u�t���x��&][5nD,.*,/+��D�i.��9�M&�5���*��Ȧ2R��V�df̙5뚯@B��A��3{�LE��ƫ�D\�	f��8�	onQe��ic5mK�)�IUU�"͙5M�b1M�%����D2�Ƣ����ήk`"C`*��$�?�(�31���Z�����-��&vq�G�(��¡P$�&߫�M��VUQ���=Q5 2����_�U�    IDAT�G"QTub�{��TXP0+�)��f���c�PA��ژM&s�f��P�8��V��A^nnjJ���C��a"�^��A'V���tff\=ޢ�L)�4��1�?�jr8S�)����_	�I�'L/�{]"�^�1�9��Z׸��G��1]g����M&3^c5<�Ֆ�JSe(E��
~d^���Led|"�e�&ćw�U5�#%U�^u��̎�TYuT�&�ʬV����e a! G��El,��?��r��9S]�2f��h4z��񆆆qjJ�LfGJ*J�I��X,����]%�L4E�x�J�	V�'d��6�]Uǳ��������������ڴ���v%n(�bR�	�;�=��h�I�H�9"M4�8����L�1����}�ر��⡡���A��Ν;�D.\x����v�3S�]�c�XKk��b���nnnF����-*1q0�&�C N��4�LE�>A��8�0�+c�\JGG�����C�-_�����l�h��w������O>��Ӯ+LPEU�fs���#�?~��p8�v�ϝ3����2W�����?�qnn��+����Z,����wR�3�SⓈk*|��O�*����%Z�TD������?����srr֭[7��T��Gy�W���?D�ѯ}�kWZ��-	��������54�3�� @�/\���?�jͱc7m~��'o�m> 8����,��n��˳Ym������u�@�f*!��-���L5��$;�����ڿqq�?��?̛7���&��~�颢�o�ۯ����߾t��+U��(�����ѩ���s��w�e2�����v��l�z�ǎ����a��Y����N�|����?�"��$&d��Q=�A��$$y�:
�"��֭[5M{�g�ΝoL(��TU]�fMuu��͛�lٲx����$dl,�i����ID999��yV���� ��Լ�� x�w�ߵg�7���LQ���s�S�`����{�./+C�7�z���n��%�������Xq��5k� ���o������**�UU�z���/��˞��={>:����{�.++;R]�a�ŋ>�裊�|����[�<��c˗-�r��Rcz�D�k-�i��������Ϸ��dgg�]�V�'??ɒ%K�,��(<�@jjj}}}WW�hv0k�ٳg+����/�������m��u�s�Ñ�� ������B��t��#G�*�b���}o�?��=== ��ӳ���~������[~���x��D����O����;�%���/�����K��p.��K��/;�������:t����F���``` ;;KJ�'�e�9�m%���^���]�akk+ ������������&���t�O\.WVV���@OOONN����j���o�����'jj�y<��>�ȃ��kO~�����{��5��Y�lS�-���5�7n�|��%��#L����S˗/��>����lC��ի�Tikk{�������Ο=���Ɲ=kVQa��^j��p���3g<x���'
]j�T^^^XP e����Ec$�'�'�޽`�e9����g�8�X,w�\q��m��w�ٺ��ͯ�:mZc��n�F����@(��z`��\nn�;=}�������h4��֎���6��v#�3��G��F?<th���P$~BD���{v��}��&?/�����_���_�I��agb��k�	wF5�???_X���������X,W�s�=�L����'���4�D"�a�\����#Ͽ�bUe�_|�+����6�@Ƙ�bѴXww�X����Ͽ�۪�i�������������:���>c�4)s�PC	 T$.Z�	��)��������������w�Y�~��+��Xl۶m˗/����cc�\i���������.�����L}��ٳ�rs#���b޵{wjJʬY�z{{C�Pwww��{���*�9s漳}�˯�������mll,�/yIc���t�\q����}[kۧ?��b�y*�HCQ�n �%4@�woI�Jp,�R���u�֩���K/���\v@,۹s�;l6���믴�sm�����UU�߷��W6���]�x��y:33�����{�mh8��?�Qss�E,�m������6�m,K5��sf�ɓ�sN�l�x��Q$��/�1�xѢ�ݶ��i�a�9���t��<�|Y��k/>��_��!'�4�NS�/Q�����|Zm�3=W�yx�������^FF��>��+V��v"ܼy����#��SO=��/}�ʉ?
���Z��4�����a�sUQ�v{<'+����(--�d2�������N��f��|CCCn��b�p�;��DqD��b1M����Ϟs8�����<"��b�ΞW��WW��pq�cz�����E� P��utɈ(
���>����ַ��F��������w��]NN��i���6��s���SO=5�eal�+�2VJ��f�(������"~��p䇌��!�K�.��v���ѩ���>p���C�QO ������'X���X�kЄ \��%܁,
Y,�+�'�������~߾}�6mjkk;��X�^�bŧ?��e˖����Ţ��<"��_�x���)�O��uKɑ��C��Ũ�?��cD����b�P(hw8�\�v���ׯ��[ZZ���E������[�y�?4%������?q�d(.**X�d��zjYJ|2���ۤ
vq ��1�
��X[�TU-)))))��J�L�v��y��ϛ'�E�z��v!2@ �"@HV�?�iC����  �F"~ߠ,P%q�qL�T g�%1�#��5-��dUS�[Q���c@�8���#s@G4���G#�֘��B��o�/���%qB�3�芤
K�@T0��β�!���V��f��>�X4
¡P��$$��e��Hb��H� Ɓs=ƘTpM���PH��f
Cd7Z��x�w�sY�[▷����D�8��4-�B�����"zJ����kZ,K,@"!q��Lo�r��@��I��8���FcQ�hI�1Ӌ���K��A9�a-�8��D�$#Q P���#!O<�^BB�`0ѥ��L�$��H�#�3H @N�Ȑ!���$!���!��!c*" N$Y&!��?�/4# ��"c�9p�[�Q	�DYf��TU4[�H��@I�����d�Ţ�m�JH		�(��L2 2�D�QY�B�&���H�� ����%i$C�S$�$nv�N���8r�i�$g	� ��R!Nz)�$���"��K�Z�}Z,ɋI 0�@�W�%��8�Vh7�NK��" c 9p4����9�ĭ��0I-�EhR	�!!��_�n%�$nm��@0   b���H�`F��P*1�[�d,�{�3@$ ��Q	zar,!q�*�dh1��"�����9u������������H$��z�~oo���Ш���Kwww8�www��PH��Ĥ� �i�h"1a'Ni.Ֆ�^۵{��=���~��z�{oי��={���o��ɓ�.]�O���盚����o������[o757K)���P�Oe� ����`js�.\�g��`0h��ϟw��eee�\������\. �#�X4�QJJ
9R������8�P(EIII�+}��|םw�&�]w�����P8����n�)���p�F���� ��N	8�h�9�UqQQ8���˷�8����qǎ�=^���[u��V�q����\�����˖Ϝ9����ܹsV�m�ٯ��F ��>�~�����tz��w��~�����ϟ��ֶa�&�<
�����ٟ�ٻ�ܹs�H���䡇2K�I$�2���T�RԳ�ٔڊ.�+#�����t8:�;f͜�{�m6۩S��}�ɒ� �����g�����կ~�j�.,,,\�rśo�e6����?������q����Gy�b����{Ǐ��3g��;g͜�rŊ����;v�����+_e��߯���iiRT$PdDzM�Y�(I%��L!L&��y�?ƐUTV��`55�::;{{��PP��JMM��l������5Mkoooll����Dy#ZU���?���6�4�RS��P[[���g�Z��������ŋ7mD�c��S�H��#�*D8��"" �)�@6}����x�n�M�1CH������_}=nݶu�l�Eq�\,x���/;���gΜ���ml<��	UUL&Swww�/nZZZ^^޳�<#��H$�X+٤{�&��X2!h�h��\.WIIqmݙ{� ,K0��>�����Q����y��񜜜%����/�ڽ��tffd������744���t�����ԝ9�3�L�Vݱ嵭=^oc�y HII�VU��-��v ̝3G�=$�y�n�R�y�%�j�1$�7f�^}�{���%Ƌ�&��SPPP^^��Z�9�������s����ɱZ,���"<h�ي�����#��={vYii{[���/,(HII��x|CCUUU�gp`���r����'///55����8��}���ԧ���q�]�]��Ԝ�l�u�I�XŪ[�������n(;�� �+�<4�_��S@�C�L�j�z������ҩiZ4�ڻ���|�	)XqĢ�Q?�H?���s?܅��!SGAx,£1%Ȑ[�Hoo��o�CC��}DJ��N�/�  �s4�%�x,���	n#+--m����h$==]�9$>f(&���Jz�8���������/1`2���
�<I�*Ék1 "d�ogU��--I��಻�ĭL�ċ� '�3��" G�����k����-�0MK��ڌ�1a$ !K��׸�f��HӴ$�Z5E���aL�J ' ��p��#B��y[�B���]��d�N�z?@@���3�*�����8i<fԯ�4��9���R���!�ȁ�6"�?	��,�/�I"��菐�pQa@��9�T8��0A*PH�#�zH�#!��E�P��"N����Db��H �8GC���ɗ���~["���L��C�$TH���$��3`��@��2�?�  0F�E �ǣ�2?CB"9~� Ś�^-g�k�q�ϟ�>z4����ݵv��(�V�U�HD�+�֍�M�-�TzԞ 8"G &�O��x���W_�RUQ�b���]Q�#G��|��~�����W6ȷ+1�n��Q%bh�@�;�O��]jj��̘?��(Ӫ��kj���m6��O�<��ӓ���`�m6������6�??k��cǎW=����|��ӵ�nw��ESSS�'?�'m6�+W����� BGGgYYi�3�S�l6ۚի,��Ĝ1}_��+�$����z��oxm붎��H$b�Y�rs��O�.l~^�����>
 ǎ۲u���p���rss�sfϚi�Z��pQQ������^|�¹s綽�z^^^gg����X,��]MM͹��7mޱsgQaaݙ��{�H�HT�������9 ��\����o��_�����ſ����i��v�333
����̙�;���/��׮Ys�ڵO���NOO+..���-��m���MM��hT�y5ǎϟ7o�ş��S�--�mmv�m�EK�,�>}��3.\�v͚��3RH$Vdz�1`��D+�S�B������ş����tmm�O-���l�088��t�3�ry�@ �⋿���p:��*6� �|hh��p��(i.�� 0�v��5 p:��&w�J$,�q����H@9Nm2U[[[8��lN��l6�Tup`0�66�Wu��)))W~QQ����H$���600�|�2wzz�^E��˭9VZ�ڂ��'�3�e�x��--��P(t��YA������ ����1���Ȇ����SYV���핍�~�ӟ���&;;kZUUUU奦��_x1;;�����_���ӧ�,�XTX�E���ADN��������
���x�b"����_~���]��q.�ĉ���^,���y�/���;v�<q�ܧ#1c��#F��U}��H'N+�k���q�5L�<�q�Ѥ�b�Kt�0�L�OL�}P�h4����E�QM�f��a�8��v,��b�h6�1����*�"F7�͚�q�M&E"Q�ل��'�	�Dj�������D&�� !1B�|�c�1��|ه�`�e��$�ɤp�TU9/��]Q�%D�X̣'!1��Hz�7Pu�	��s��1	��/C# ���Q�{[$$z4#U������#��H0�zS�DJ0G]�!��$$��3 P���aN (wiJH$�)1�[@��	8ILB"q�L�n1��f-HH2�!!�O�eB���%T���D�X�s�H/�#��K~IH$�/��)qi.JH$I�!�z�z);\�*��H�"Ӊ�青D]S��H
��ؿ�r@�+/�`2�!!�CQ�!m�d�	�dh2� �1ԃ�dt��Y�;c"I�H�A3$NH�[���D,E�P9� PS\�����ع���l8�dz���/�|�P(�����?�ʆw�u�]�����"�.%nb����H��ŸE�c��2���ojj��h��{{{M&өӵm�mO=���a���{3=���sw��#_��Mm-[YT2T'���c�`0�q"��ZXP��ݳo߾������=wݵ}��������|�f�mظ)vtt�&ӣ�|����hM;���A�_���<�:u��]���TUU>���?������O���o�o<��R($��@��g��E�?QhqjY6s�L����_�ǫ[^kii�x2W�\y�k���3����7���6���� ������}�/J��w����z�}o��=�'O<���b� �������~����ӧk[[ZfΜq�S�`���G�iN�SʄD�ME�ĘأIH����)_s��?���O>���o�?���+�'�XO�w��5������R��9�g������)NgEyy^^^�{X5�L�ں�]�w�|������LwzzSS�������du{�I��##;4!ޱe�W��6[Ue��y����L}= �Bt�N�޽{�+W�^�����S�*jH�p$��F�)���eːoh��u�f�$"D�5{Vùs��g�̝#BbRb��cz^��䳩������hkk������())q:---�`0Gc����p$r�w=������5�/\���4,c
��}}-���Ò��ӵ�V�5=--����~mm �����曱X������===RX$��C �y!�\�+!���Sk,�춖��Nq:>��O���9[�i��~�����-������@ii��	�geeeFFƳO����SU �M& 0���~��w����Xx�mi�i ���WQ^6g�Q�$�FcQ �bZ$�D#ш�eKQ��#��.�6 @�A���f��6e��'���?}����o��j���D21�:������N0���� ��p��+�b��'N���Ι3f�Ͳ���Tyc̨����$�D��q�u�3�\�����9�g]�wBB�Fي������(��n�=d���ʊ��
��%�\��0 D��i�F�i�	k2 DBH����	L,���KE#}0bR�IH$h*�I L,�ʋdS	���z���D�`ђL�H�&�:�T���.$��IH$�5�ܢW- 2B�A	����!"�Ԋ������^;Q/m/��" 7򩈒\�#�D�a��%n�l��d���	H��P��Ԩb�����oN�VANNNR8Fz��P%$  FF��d�c��������I|��0#�A(ve"!#��,�hBBB"1k�!�e��3I�IF%$�ƐHzT�4@$��'�>&!����9 q"b(j{��z�d��DRt�^'PՌ6�`�cL&,JH$l.2��b�4���R�IH$�\��e���H���,�$!��O���1��������Djl��//'��D���$$��MG $�IH$A��ȥU��D�`"�CSB"9�Lwʀ�{�H��0��P���><���D�e�m�I�/��� #D�> �� �����o����&{��s����Oʂ����2�o�    IDAT�� �C��������omme�RZRb�Zc�XSS��aw��\�������2�JJJ���:;:���(55U�$���� ��K�
��kk�Μ����)+-�U�%�m'�7i"$B�C4r��(��z7m��ѩ�۷�ܺmUW���뵵u����<��׷i�暚c|���������>u�tmힽ{���+q�s```�ƍ�@ >��P�������5-&�Bb2�1 @ �#1=��@����'>���Ly��τB���Ǎ��o߹��_�bvv���D#gc�?�(���9D\�l����������������_yZ��^YY�i�+WHq��s��
�*���A�Qv%T���'+�c2�L&�'�����ssrc�%�x��n�ժic�s~��A����p @4��*!qCi�H�G �zn��Zp�9�D�r�555G"�`0����+�r��I�4a�������H$�9ܽg�ի֮Y=��:2���@4�4 ��
q�X,644$B���!q������"}JE .B��@�0�����������Pe�ŧkO��qS8�=kfii�]k׾��+���N��m��������_�`�Z�l6[vV֦ͯ�����a��f�x<�mݚ�����������~��w�j����x���h�w�mhؾc������`�7Ͽ�أ�Ia��.%�w�U�2��$"��sL��Wo?9s���h�e6�23=��e��ӧMw:eee,P%??/??/-=M�i.�k��YU��.WjNNΙ3����i���\E��K�.���%PTU-//OOO/**Z�t���III)).IIM�x<99����v��j���nUU��򲳳M&r�Fk[[_��Ǆ�Z��M�����������m1��3�O�IF�;#��g,���f�<���9s8猱���ں���B���v����W�mt���?^����D����8�)N' 0�JKK�HI$�� �����V�
455��m��(���p��]��5�m���W�[������R� �#q�Hp�gWVV��7�!�?a��_��s����"߮�M�1yS t[q�����[cf�y�'I):)!�DC�G0���^��ᔧKH����P���#��@��LB"QEf�y&"6��/��IH$�� ��� �%��� ��D�l8��p`���*,�1	�D�h ���"׷Es�x�?		�D��p��z�{���P����H
� TBѲV7!���cI�	 !r���#pW��H�K�@�	���pDb �d�?	��5�0IE��"r$M��rǰ�D����qE���4AZ��ۉ_	cF���$	�K�IH$ �����DM��}d�6o>y�#�{,۰qc{{�o�u���w��8~�ĕ_ٻ���cǓu^�����rk[�+6�����9������4I�j+
L�vכI��P5up��>�� ���{��|ZZZyYYffFII�'�s�W:����z�u6�mƌ�N�sڴiV�e�����1Y�Q�ʐG��)�o\���5�UU�G������'���9c��bi<�x��\��}�}�����;v�v�����w�飯��k����ԘL��z���P|�?0�}����֊��;׮u:����F���g333|���Gk<Y�ٳf���:|xႅuugv��=c���Ӫ `���D����������r:��/\x�]����щ�'���@���w�9s�̡�����FC���>�����]����
e��'�dH�{����2����V�x<V����3�=V�r�팱��§�|2%Źi�f"�x<[�n;v�x������B�0�2��?�ؼ�s����&U�3{��=~���}��.���?���p��7�t8����b��A�ż`�m�~�'N�����������z���m��=�mm6nZ�l٢Em6�g>�~��;~����^o$yg��j�s�����/N�6�εk���fWw��O��H�y]F���F=l6[YYٙ���--N�3## 
���5����w�G�xo|ߗ2�ľ � wR\D����Z����m{��s�0�4g��m��������������3�����UU�HJ� ��D�K��C��e�"�L *Qb�$Jd�E�]�����lme�9��9��o�y���^Us� ���wzzzeu�X,aR4��O��m{euE>x�������}vcc����P,nll,,,�����G#���1�uWVV�1v�ĉ���K/�R�������'��9s��� �^\Z���sG-���y���Z[[3��ݑ����>����|�P�'�����uDQ�8y.ѷ9�ϝ;{otl����'�P(��?�y4�p�|�.F�P���#��$����R���B�K/��דߡ3>1���u�>}�4��� ���4��ͯ�����߼�����'�6�.�Q�TB9�  \��?������u�����6$����a��������?�������n}��!CB $S�H�<��G$������n �y���0 le2�l���p�T�m�&��05�ҋ/~x�#!�i������WV���b)x�յ5�0:::��\~²�����ׯ��������X4��ڒ��%(C �Ύ�������奥\.W�����>Ӵ
���R8�������D".G���O?�\�W�w�ރSD�J��^�F�s���'��"C�	��BH��o��1ƞ��D"��� m���G���?����]����]�~���_���2����⹳g�/,<�����_��7������s|h��������zcc�4\�pX�j��zD:6��H?���x���F�/��/����VJ$rJO(������/�����_��o��ڒH$~��7���������ʹL�X}C3�4h���'��������y�=�T*
W�]��� 02z�������]��9�_��*��7z�7BA��s��.$.��yW������3t5�6\�������?��Q���!��d�&�"FRdТ:K�i���B�*}5�ͯ��HeYUB��l��x��9�d۪B���lz��	d@VU�����k<Up]�q���1�m,�d�I�3�>뱞Z׋��T�P,��ՙ��� ;H�[��m�Ӯ��u�xz��dJ�R�?��W�ӷ�Cj>UU�b6�K��z�5����\�w��2EV~�K�d�RiiyI��j<=Flu����o& L  �P�Ū'H�֙����ML�R$$7C� AF58��bi��=O7Pi|߽ĥ����Z�$9Z��2hjN� ���lai�'UC�۶G��t!�(�	٘Ijb`m���޾;����wB�{�b��ō;O�x�c"��b  �� ��C���~�[�o��C��׽}wdiy�v�2��`��v]V*��j3���W���@�5�71����g�>5=��S-G)��^0�H��i��b��[�\���@<כ���ٹ�{�c��[��5ȹT`
A�	ɏ������OL��/=����E5��w�ȱ�����Skkk��8���^�3�@B�,�
�oo�RP>��y����d{[[SSc}}}],
���#�4�4p!<�-�J�\nc#���X[_?�fY���d=&�c�`*��������lȲL�d��<�QC��@Bp�]�s]��n����`"��!��(��΂h<�@ "D@ d�`�Ld��hh��>*Q���*���Ye�����ޅL�b��1�)k544��'�"� � rD0	b:����_Sm� �K�#|�ڎih��S$��I�<P j�Z��2ɋ� 2_���e�&�v54��+J�P0��	��4�}{�H@D`�Kh@!M�n���ؿ�!2F�L%�_ ����_+�1e��ɜ���B��q �FD �RQ��ihh�X�c�C9σ3��c�,�4�	  ��l2�t�^Cc߆���`�=5I��1�}Fb�9���{���t'����Y3$PP�&q0m�Z�Ta�,�@٣	��Gm�44��,�	o& !��&Y��˩44��!��HL� ������q ��,�b��?s ��#ihh��Wy�Lh�_	��B�����ط)��"�2)h����~���$�2
#$DyqF@��KED�\.�H8���_f�����z�w��8�w��][]�B477�:u���7�����Fc���I����y���޽{筷�����7o^�tQ/�ΰm���k����������̱���_=��%���1DQN��Y{����*���}���\���۷n߾x��������l�o޼��_<B������'�~�馾�����!����cXs<&�������/�����5 ��b/��³�>
���L6;|cXrjs�xhU����*}5'(��xL��3 �Sf���ﾷ����BpΥ�,k;�"���M�q�T�Z2K3����BҰACH�=��5>>	�u��[�E��Db�!1*IC2)���j�O��R�T�#~x�ƍ��uuu��������r���wm�)��έglWP�~�	,$�  ���E���oB��ɘ��E&{���&�e��<r�왞�n�{�4�{.C�k2&׼�ӎ1f}��
_�4M���mٱhd�	'T��H`
H��A�EȢ��o�111���T( �0�d2��ֶ��`?9"zJö���_���|� ' �,��'zz{����l�O��)�3�����k}=�0Ξ={�̙���?� FFF����x㍾��j�쩍7Z[���ܹa��U�������v�;'�~�3L�P�E����Ν{��C!�ҥ�--������^����^z���#�a<�1�����_]_C7��4 ����1�@���3�5�G7�1���QWW���r�P��zjyy�ĉz�w@$�����v��."&��ӧO��/777���ΡT��6� &#ÔY{"&+�h�^	3��Ç �H��G?�L�hl�D"q��˧Ϝv�,ˬ��3MS��wD�� Mٜ)˂�Ɂ9���F�Ѩ.�6�M$z�?!�J����	2"��15���nM �%AZ�44�W���
@�����q`2*w/;��1QN����_!c�B�,�"=5GC� 2�cdj� ��#���ih�ێɎ0}�?A@%�Tp�EG�xkh��! ��(�8�y;�xEA��54��*JN	D2��/[�BxD��O�<44�k�0Uw�e�=^����1��2"��b���]G�3����C�(�6�p�`��C� "�L���>���k7�C�$�r�ޅm�-b!LD0>�]@T�L�'R�Y��g�u8�.y�)�.P�!��3Qw�]��ZPeݍƉv#;�=v9<X��k|� r69q�i�v��a4�0j4��-	v0�F`I0��*���]���o�{����J�#ۃ�"���ק��!�L���cv��hb�1�B�]�֯��S��"-n�/g�c�ƅ�5��!j(SU�Ws��Z䱑�Oyc+���}�<p9Ϲsi��`�pS�b�-ѵi��w�ކ��4��-o����ƞ�䉀�Ą��-�E�cc�JF��sO��Ե�xwľ�P��LI��}k��v ��Q�;�g�=�'ʩ��!�{���ȋƜ՜��}<�N�x�F��[�?<H�\�6��Y�{�Q�y# �)�H j2eE�>�r�2:�q�(���}w-���r_̸S�zj�����괻�)j�/�=�"�!��ܪ�����k||�k��a=/���o��]��<�!~C������w�F1S<��3���F�=��}kB�D��i���b��5���i�]�s�Fn���.G��i1�Q�)C�WД��.���ߪ|��U�.���':Co��Y���o����{�č�:6��
�w^c�ì�ޘNy�� �G��C�mg�Υ��V�^��l|��?�(e�ڽ�.������ZSw`H�&��"$"�U󮰰��*67l�囯�6���C�����/f�减��ސ��#�N��M�x8�����#k9~oi/�����P����� y�Vo�u:v}��r��U�7Eѡ��@�RF�fh�c�͐����ǈ���2%qo�]�� �G'����k�7=��,{��!�|t{�q�p��F�����
�3<oS]U ���ja�J�$!"��ry��rU�$W��  �62���j�Aw��)���p��(lA���ljw��T� ���l�{[AhK�]I���Τ��S�G"�EB��gѥ�J�G���gt��Xkש��n[��'�뒱�x��ͨ��^g���]��L���1���Z������կC_��?����2 ��`��ĺ�\�l�J��_�K& !1�|T�-m�r6Uw��w��>�jξ5�<�g�yּ��Vc]��g���|O�� �l�2E�g%�Z�l#ω����E-�G0�Em	㕡H�D����K�:C��杣mV}��.:�7
�-��
t{��E,<s(���8�=��cVG��.𻋮 za "��Yw���rAóv,��{öKW�v�f\�V���	��*q�;|�պ2^d�..�2p�
�TNܘqr6�}:Zy�#���З3"���^p2Eq�#�^ol�Ȣ;�j6ֱ��pc֎Xx�#�cK�����;�j�7���޲��[�0�:�:e "��
�#l6��_{�&s��:}�>k�I��&D2�a����Ҏ.J[�a�ۘ�r �*
NЙT�9׳��#�Z�J��[v��Y4�B�z,�	�����l��)�D���1�r6��2�ؕ�RO�2�y����h0���+^p�l�Yt����ڱhW�XH��8[���LO�̡�t�;��Xxc֩xV���ز{z�>�_�=z�/l����v��	�Kj����צ언���X��#m�b��7R�.�>�h�v,ҕ4��	~4�N
�,��dWh:��Y��B�)�bo8l�JFx�
6em��<m��TN�q,��_��z��{Cs���H[����R�!!`� \� �&��F3j�`��)���u�+ՖZ�e�&��+T��@��zE"�Y������� �2}e����qf9��"Υ�_�.z�"]h����Ж0r�h����O�D<̂�4��~<Y��G���~��؏�Ō���?;k�7����qs���	b�F,��b"� "��z�2�����ƁȘ���g�������;���z��!�*��#>�,��g�Ap��Ai�����rb��<�f�[z������ AD ����E7o�lڛXq���Ѽ2^�\�^;9�����[���'�K��^�|� 6���W�N�(�'ཻ�D��l,cO�������04՘ ��ǪUD`;ء�t-�l_�X�����*�H�������t~���x�q�|�h$5�g��v2�Lt=r8Qŕ9���=
���	O�푁*StH>.�N 9[̧����B�N�g9��B�����"��r��n�#�.�f�ݎb<�^��Cx�h$��j��>����� �;�b2F$S��B�l��2#I�Bp9"�#D�4��x���b��A�vQ<��<֞�}&��	Xy\p��� b����	��1��C�f���,_��Qa!���i��ݚ���Ӷ���:CGZ�dq�h0�:���|�sAW�&̓����ǿY�$�.��ۭ�z&s�+[<5L2E�ݰ_<���bھ6e�p�h l�Zf �U�uv�p8���)]�XuC&��l�1�x��㡤��b�ø��R��"1�C��+bbɥ北�1�_(N`�ԙ4[F�(<A'�B�;C-�L�+8����;�c��C��-^rI���V�|bof���*eL]?�:�-bab�<�CсV+l�OƂN����4�����#��<\N��I���K����8;��,O@��ܷ{��#��F^H��KB���KW�J\�蒛�ť�P�!��	D�r�v��R]/���vI���)��#���a��|�Y��پ���Ѝ��n�{��vMe�@���J>  IDAT��s����O��D1���C�x��ڕ4~t*z�px:�ݞw `d��i2�a6<k���q�)	.�Ƭ=��_�UǸ�[Nc���		�+c�x/��7��Y�����Rɥ�D�'�%ۥ��\u/�z�M!���%9=�e+-u5�V�����3*��#�s��^}{`מY���Ɲ;��e�ϯ7R�����] �_�(ܕU�}_1�j�u:vu�ts���~,c��Rx����S�gSn�.���fC�bc����+�J��6��z)R����F�_���"2��΀eD#ӍX��6�N;�{�������S��-��[�j ��,��C�:XԪV�n���y��Z�jGW���W&������5Ml3���lѿ�<��V��~���=�"�|��S��ܡ���z�Fw�_�j������FM�x��:8 �  2VN�߲���2��c��y��$g �����6�)�;;�{�-� ���4�C�j+P�5��{b�h[�k�>�j��0�.��fЖ`�z��ni��v�����|�ߪqjXE^�P�̽j���:l��>�P��w���KVS�,���^�h��=xD,|��j��Q�Q������%�5�O4���!���ikv�h�⫃���j�W<��Z�M��f��^�NvԮ���3P��jB01��;��8{�T�T���<�����u2|��6'<ƷO����ݷԨfZ��c�g�k(�xD�T�L HL 1 �U��ݚ�2h�׳�9o�(���=@6���6Ov��{�d�Vg�b�]�	O�v�4�d�q��l�c{dG'٤I�`T��@"�{�e�X�|��x�"�y�J�BBo��;21�d�u'��v�!�/+2�X�q�ŘJ��k|� �%*�9�z����X֝4��XS|_��@` �&"� D@��ߍ�8�ek�lI\�S�5v�IBDCc�Wɻ�4`���o1�6�l��.��Q�BXw�����& &d�������:֤w�[�ɠ!��4�{�c�@�b�g�t��2��o ��r{C�h�1��2e�P����{`r�����Dd P�ET.�H�444�i�ԕ�)���gD�;����FY�P�b��"�? ���jh�G�*�`JD�Q�J�}�S;�;���_��Q�v��3����e@]�a�eh�RF������+���}BHo��QQzw��1_!C9}�P|Ы<]y��t]Վ2����B��ho�?tPjO&HR	$|�}��R��Dծ���� `�1��.H>��3^��Yk���|�[��Yo�ݸ�c���yo hJ
h9bQ�%�MB�@ABk��BB�؋�eKtu��|��to�[�tpь� �>�&�_���恩U�3���"S���,g4]���-$t�6���V��B���	*��X����[�7�ɂ��Y�2%�`�]�|����AC��) F|׺GB���F�ƪ�p}�}�����]��������Y $�k��t��:����]��<m��!��|���5�/�$���q`������U���o\�vs\7���f!Öb�ֵ<5a>-fӵu��>�U�� ��U�,���Q6�Mm�J��a���������X�$f�_��4_ڍ���8�h�c�����Yt&W\�VXD0z�L���&C "��w"�r�j�;�Q��-�z�j w9����7v������M۶�a444��_�|9~�D���d�Y�X}}�ɓ'��������������fe9�w���s��~��v-G�`ik>��z����f�y��d�H������󷣅G���#"�1kKR戅��¹��9�i����ó��G#�=�%Ut�#�֑6���I"U9l�پ0|1m��dti˓����R�|��"�3<gS��.i��� Bne�S�h�L��yW�^�r壖�ֿ���x�ȑ?��?vl||�׿�u!_x��gggbG{����~�k���������0�@��k����vT�m������Nw�Qr&v�YqN�\q{�����{#šv�r_��;֮���@��A)�&�r_��� ��C��m��`2�������s�׏G*��:��z 6�`Sަ\I|Wn�ٍj���/D 0���V}E�s�����W��:u��s�=����G/={���巿����ȅ���i��p�"޺}��\��7�NoF������Ƥ:�\������P_���C�|~tt���.�J���?~ ���f�g�����]]]�tzrr���ѣG��Z'&&��<� �z05U,���O�<����GG����t:����$$?{%�+��������_q;�Ʊ�нw�a�ڈ���fR ��
�ֲ�%�.�W����8�i�C&R� �;B�ul=������F���q�%��d���W\�#D�m2Z�t�ׅ�Ȣ�.���1�n�V��'��'���E� P�y�A�b탂w|Ǒ��d2�̹s!��<OZ6�X������D>��)SSSW�|42:��ݍ�������߿r�mہ^Z^�g2��}����r�X�v����x*����///�����{?�˙��9��r���fzskk�w�qgii���`j���V&�q]��իwGF��������lnn>1�6�v7>�m�!�ݚs��Fc�Q	\���FG���`$�ly�K=��P�Bo�2�C���p(i�~<z�Ք� ���|i0�)�͢p<*9��5�i�i2 �+i��d4e�-�ۧc��[g�C�0K��O�Ē1�T���l�	ܙ��Z]��)*Ict`��KK���X FGG`|l�s��}�}�m?J4l�f4min���]�_Yօ����ʊT `��9s���%�А�e���  ����K���j,[_O�/T��h4��Ҳ���N��!"�f��l �Ɇ���'�.]���9r�H<^g����R6�][[{�g^{�����'B�p[7r��nl�YW9[��ο���K[������5W
I<�7�7f��G
���!��6����Y�>m��^ˊ�Eg5�7�b5��.�_����FNd��9n�¬��t9��N����L�t��uLҒ4DY"�DL?���Z�+��MD��-�3��aHo0�N3ƶ����k�kk��+瞞�˗�}�/����������ٶ���]s�%�ʇW{�2f�$D@d!+d��<V���~���6<|���k�㚆���v�������z 0M+
	!n߾}�ڵ�����.�뺌�H8,��I�c�������2����Ȋ�u��Y�M�W�B&"J�S�����8�W@�A4�;Sfׅ�ۧ���Ny�&LB�!�2�<z������������Q�1�1�#�S�J466��i��]�t����7��|n}m-�HX���S2��������^�1����b$.��1�\�Y^YNo�C���D�_}�q��tOOOssS.�K6&����2M���Y��鍴d�q �z�4ݿ�`}}�I�c;PEKL�>>gg0<�N�y��\�z7g�kSv�wD�%Qt�dg�X�u�ݚIy_ww\.>�o�ƍ��!D(��7��e?��GXG�Qa�Gr�� X��q�3t�Ք��\@2�\NR���M������%�.�пz&��D����[=������ ����?�\��^D,�J�����cu�ʟ�BSSS|���;wN�<y�ȑ��֎���w�lmn&�ID��:��fg���fffFGGZ[ۤ��!"�,�0�.���~������ӧZZZ^��R��~����	2MӲ, 0��ѣ$����XԲ�p8���omm���455���o_�p[>蝧vϦ����L�<s(4�n�]p2��#���}{x�!�����裉�i��G"�9qu�D �P;�~%��S�Ȣs��j�w����p��c+n]�bl&��z�̵D��Ȳ��@X
$l��cŎ�աȉ�	�1���u=��� �w�3���J��ٖ72d�����|��R���+�L���T��ի�<x������
O=���F�0��ە�5a�q<��b!�fA\�*��X]I�ּse��De·ڭ��F��B*���^V���3S����` 04	Dy�) ���<aTAV�� �]�H$�ҋ/��y5��ǱcC�Z�j3b��l�]�>������)���[Mu����B�{�Naz�{B,a'�B�cV*/��Ob�^�|���T&3Q�l"1"( �u��#U�C��Ut"�H$�<�L&���f�v̻T��UO?�,)�'�|	�n4fֽ/gm�ɻ��x�j>�ՕMu�,��7�Η�T��k�<Q�`H����Cܹ!Z�A�_߽,���@�����'yzYWu|Ј���QN!� `�
�I�A�l���*V٩Yk��F�^"V��]Iv�W�As�,�8P-�]�6!�*0&k�C�@(���f��s�3�Ecg/�ʩ�|�9����D,|��jKT��py1](ؠ�i�0$B$���!���l���X�QШł�Q���!�p��>Hԅ��D�|�D4�`�T�+Ǌ2��ф� �Kn���L:;�`��FDfh�� ]DfX�zօ𭓚��t��>Wt!�LM�p+�?�%q�q[�%N.�@ �X�P[�����W���į��3���L�J-u,S��Kz�� كO2_9ju7��1��s�}tOpd�:L !<Wx%\]N#
����ٞ��ڨ0c��1:��pװ= p s�C�-�t�Oj>��*���i4[��M�^ul!p@ M��B�@��  !�gK�_�u�5ּ3�V̻=�{g;�̻78�f��|��2�����:�u��l"�N��M���_\O&p�J:5(����C������6�Ay;�8�H���C.k_��;v�+�o�$F �@ )��V\��D>c������;�3s�k�QA�&����m�H��4Q����V�uE�@+ө*�m<��������x�j��lϔ2������*S�HL��������0NCC���Z����U�C���E9(�h��|u�r�) !����YWmnM�{f����g�_����Ԛ��B߈I_�h�Ȇhd~F��� �͗�Ru�h[g�^Y)b��w~yc�������R�\� h4G�5���L=M%G�[�MEb���zƴ9�xڱ���������"���8�� (�$2��G+{ 	"[�D��	�l�OO,�vgws(��O5�Rp���.��/>_�� �Ƃa8��&ukŌ��1�y�dk4��q�LB
D?�!��Rfce+^mh��)���;D�K��������f� T!���X��h��'��	��IV�
U������S��w%M�i�1��|岥�[sW?M���H� Hva���(g��_�C?!�G '��d�
:�a�|N�!Q>r��ؙ�d>������p!��z�έ��K�V�K:gd����a`f�<��2�S�y%|j$$��(��"�L� $���!�K$��ǻz�[���PذB�a0�@�����@p��p]�8^!o�Ϧ&F�6�%G�'�Q�jD�\��	uM 8��	���*!G��y~M/"r9�[ A@(䅵 b@�,���b��X$j�,��J�����VS�P]x���B/mnE�L0�����d��x�zV�B� T����˴)����#�X�?�*��uS���g_�<���ݒZ�G�D�Hm����{#<�@E�/V~��|��T.�����~�[�O=\�_��F���9�D���CP޲��8 	�( "Wl���B`��&c��+^Vl?F���mA���q߁�.wl��ۙtas3�:��(2���k�d8%_�!2T<  dʭ�`���B�Lp�Ȕk��>p�O$$�I6�Y0P��+U
3W�L�������8"U�L� be�4T5�~	30�����?v��!%�����D����}h��{	��&�O  (��!M(���X�\�!F�!�*�>1U��O
���U���o%�P�CU�2�,+���6��]��`��rO�_]$y�Hnu��(��^"�l[���G pBAQQ~R�I�!1@@4X�#�?H��!�X��JSe�K.$AY��ڇ�m@�4T��)�,�@��:9��p~�;%h�"$4U���R�P6�A�ϧ������(P2L���W>�\m����'" J[�4(��B��
�cHH(@vm#C!�;Sc��I�FLZZIQC��q ��5��j���B� ɪ�Q�)�T�p�)H�1D�&J���P�a�P������A�t �H ���OXg%9R����0���S�$�\�22`�/� ԗG$ ����(��`�4����!S�R6Ի�9��`Rc��#��o��
ˍ���'�:��,�܉�(��IaF9!J���4,;9��a�U!���G�6����'_p �8�����ߎ�c�gMP� �JQ1�)H @�n؂�M�J�=	d*���gH "I�א�!�i#�҈LM��}X��1y*�Y`��˟�P����% �u5��Wm>R�*�=|�Pn9�B�o�r�Q�IR�'u-b`�P�䲋�#������ˆC���`@~]����3��|��Z��WY�W��n$Ç�v��H��_��LAK-f �@&�P%z� ��@���Azܷ���	����Ɂ ��cϤ�PPi� ʢ��TC� *�T�ک`S�?���~T�G֗զ\:��+m��Ai2�ғ	��_0�~��A(ۄ���t�-�9d0u�*}3_��7ဂ�n. S���[� C ʒ(�T��2�R/�R��s@C� �" � ��/��� �u$�7H$}�<�$�VZfo}/�R���#]��P;.m/127�B�1"(V�e$ C.-I[-?��*JF@b$��`��(#��C@�H@�����������P	ƈ��

_�SyB?R̂�Ay$!����)o%r~O�$ ��Aҟ��� ��)ŉ�U�����ȷQT�C����FE�����%�����w[�����T� �`�CE�q�R��.��}����O��� f$JjR�٪������kV�*�-S��� ×�~B@0�Uݷ��j@�M��
BcߏU2)��y圪G�� �sKR�'��D 1_�	% ~$CA�@E8( � f-�	���R��T�7�gK'�|�Q� Q�B9�S��j�2�2l��寨�Xd��H�v��D�K��_�k�/�k\���V) y�}u�G^���x9n�L�@E���ؤX�����o|�?P��Ug���f_nE��oW(~^~��    IEND�B`�