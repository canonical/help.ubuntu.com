<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Redigera en trådlös anslutning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Redigera en trådlös anslutning</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">This topic describes all of the options that are available when you edit
a wireless network connection. To edit a connection, click the
<span class="gui">network menu</span> in the menu bar and select <span class="gui">Edit Connections</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Most networks will work fine if you leave these settings at their defaults, so you probably don't need to change any of them. Many of the options here are provided to give you greater control over more advanced networks.</p></div></div></div></div>
</div>
<div id="available" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Available to all users / Connect automatically</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Connect automatically</span></dt>
<dd class="terms">
<p class="p">Check this option if you would like the computer to try to connect to this wireless network whenever it is in range.</p>
<p class="p">If several networks which are set to connect automatically are in range, the computer will connect to the first one shown in the <span class="gui">Wireless</span> tab in the <span class="gui">Network Connections</span> window. It won't disconnect from one available network to connect to a different one that has just come in range.</p>
</dd>
<dt class="terms"><span class="gui">Available to all users</span></dt>
<dd class="terms">
<p class="p">Check this if you would like all of the users on the computer to have access to this wireless network. If the network has a <span class="link"><a href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?">WEP/WPA password</a></span> and you have checked this option, you will only need to enter the password once. All of the other users on your computer will be able to connect to the network without having to know the password themselves.</p>
<p class="p">If this is checked, you need to be an <span class="link"><a href="user-admin-explain.html" title="How do administrative privileges work?">administrator</a></span> to change any of the settings for this network. You may be asked to enter your admin password.</p>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div id="wireless" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Wireless</span></h2></div>
<div class="region">
<div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">SSID</span></dt>
<dd class="terms"><p class="p">This is the name of the wireless network you are connecting to, otherwise known as the <span class="em">Service Set Identifier</span>. Don't change this unless you have changed the name of the wireless network (for example, by changing the settings of your wireless router or base station).</p></dd>
<dt class="terms"><span class="gui">Mode</span></dt>
<dd class="terms">
<p class="p">Use this to specify whether you are connecting to an <span class="gui">Infrastructure</span> network (one where computers wirelessly connect to a central base station or router) or an <span class="gui">Ad-hoc</span> network (where there is no base station, and the computers in the network connect to one another). Most networks are infrastructure ones; you may wish to <span class="link"><a href="net-wireless-adhoc.html" title="Create a wireless hotspot">set-up your own ad-hoc network</a></span> though.</p>
<p class="p">If you choose <span class="gui">Ad-hoc</span>, you will see two other options, <span class="gui">Band</span> and <span class="gui">Channel</span>. These determine which wireless frequency band the ad-hoc wireless network will operate on. Some computers are only able to work on certain bands (for example, only <span class="gui">A</span> or only <span class="gui">B/G</span>), so you might want to pick a band that all of the computers in the ad-hoc network can use. In busy places, there might be several wireless networks sharing the same channel; this might slow-down your connection, so you can change which channel you are using too.</p>
</dd>
<dt class="terms"><span class="gui">BSSID</span></dt>
<dd class="terms"><p class="p">This is the <span class="em">Basic Service Set Identifier</span>. The SSID (see above) is the name of the network which humans are intended to read; the BSSID is a name which the computer understands (it's a string of letters and numbers that is supposed to be unique to the wireless network). If a <span class="link"><a href="net-wireless-hidden.html" title="Connect to a hidden wireless network">network is hidden</a></span>, it will not have an SSID but it will have a BSSID.</p></dd>
<dt class="terms"><span class="gui">Device MAC address</span></dt>
<dd class="terms">
<p class="p">A <span class="link"><a href="net-macaddress.html" title="What is a MAC address?">MAC address</a></span> is a code which identifies a piece of network hardware (for example, a wireless card, an Ethernet network card or a router). Every device that you can connect to a network has a unique MAC address which was given to it in the factory.</p>
<p class="p">This option can be used to change the MAC address of your network card.</p>
</dd>
<dt class="terms"><span class="gui">Cloned MAC address</span></dt>
<dd class="terms"><p class="p">Your network hardware (wireless card) can pretend to have a different MAC address. This is useful if you have a device or service which will only communicate with a certain MAC address (for example, a cable broadband modem). If you put that MAC address into the <span class="gui">cloned MAC address</span> box, the device/service will think that your computer has the cloned MAC address rather than its real one.</p></dd>
<dt class="terms"><span class="gui">MTU</span></dt>
<dd class="terms"><p class="p">This setting changes the <span class="em">Maximum Transmission Unit</span>, which is the maximum size of a chunk of data that can be sent over the network. When files are sent over a network, data is broken up into small chunks (or packets). The optimal MTU for your network will depend on how likely it is for packets to be lost (due to a noisy connection) and how fast the connection is. In general, you should not need to change this setting.</p></dd>
</dl></div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless-hidden.html" title="Connect to a hidden wireless network">Connect to a hidden wireless network</a><span class="desc"> — Click the <span class="gui">network menu</span> on the menu bar and select <span class="gui">Connect to Hidden Wireless Network</span>.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="security" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Trådlös säkerhet</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Security</span></dt>
<dd class="terms">
<p class="p">This defines what sort of <span class="em">encryption</span> your wireless network uses. Encrypted connections help protect your wireless connection from being intercepted, so other people can't "listen in" and see what websites you're visiting and so on.</p>
<p class="p">Some types of encryption are stronger than others, but may not be supported by older wireless networking equipment. You'll normally need to type a password for the connection; more sophisticated types of security may also require a username and a digital "certificate". See <span class="link"><a href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?">What do WEP and WPA mean?</a></span> for more information on popular types of wireless encryption.</p>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div id="ipv4" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">IPv4 Settings</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Use this tab to define information like the IP address of your computer and which DNS servers it should use. Change the <span class="gui">Method</span> to see different ways of getting/setting that information.</p>
<p class="p">Följande metoder finns tillgängliga:</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Automatic (DHCP)</span></dt>
<dd class="terms"><p class="p">Get information like the IP address and DNS server to use from a <span class="em">DHCP server</span>. A DHCP server is a computer (or other device, like a router) connected to the network which decides which network settings your computer should have - when you first connect to the network, you will automatically be assigned the correct settings. Most networks use DHCP.</p></dd>
<dt class="terms"><span class="gui">Automatic (DHCP) addresses only</span></dt>
<dd class="terms"><p class="p">If you choose this setting, your computer will get its IP address from a DHCP server, but you will have to manually define other details (like which DNS server to use).</p></dd>
<dt class="terms"><span class="gui">Manual</span></dt>
<dd class="terms"><p class="p">Choose this option if you would like to define all of the network settings yourself, including which IP address the computer should use.</p></dd>
<dt class="terms"><span class="gui">Link-Local Only</span></dt>
<dd class="terms"><p class="p"><span class="em">Link-Local</span> is a way of connecting computers together on a network without requiring a DHCP server or manually defining IP addresses and other information. If you connect to a Link-Local network, the computers on the network will decide amongst themselves which IP addresses to use and so on. This is useful if you want to temporarily connect a few computers together so they communicate with each other.</p></dd>
<dt class="terms"><span class="gui">Disabled</span></dt>
<dd class="terms"><p class="p">This option will disable the network connection and prevent you from connecting to it. Note that <span class="gui">IPv4</span> and <span class="gui">IPv6</span> are treated as separate connections even though they are for the same network card. If you have one enabled, you may wish to set the other to disabled.</p></dd>
</dl></div></div></div>
</div></div>
</div></div>
<div id="ipv6" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">IPv6 Settings</span></h2></div>
<div class="region"><div class="contents"><p class="p">This is similar to the <span class="gui">IPv4</span> tab except it deals with the newer IPv6 standard. Very modern networks use IPv6, but IPv4 is still more popular at the moment.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a><span class="desc"> — 
      <span class="link"><a href="net-wireless-connect.html" title="Connect to a wireless network">Connect to wifi</a></span>,
      <span class="link"><a href="net-wireless-hidden.html" title="Connect to a hidden wireless network">Hidden networks</a></span>,
      <span class="link"><a href="net-wireless-edit-connection.html" title="Redigera en trådlös anslutning">Edit connection settings</a></span>,
      <span class="link"><a href="net-wireless-disconnecting.html" title="Why does my wireless network keep disconnecting?">Disconnecting</a></span>…
    </span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
