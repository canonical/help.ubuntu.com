<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Öppna program för enheter eller skivor</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#removable" title="Flyttbara enheter och externa diskar">Flyttbara enheter och externa diskar</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#photos" title="Foton och digitalkameror">Foton</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#videos" title="Videor och videokameror">Videor</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Öppna program för enheter eller skivor</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan göra så att ett program startas automatiskt när du ansluter en enhet eller matar in en skiva eller ett mediakort. Du kanske till exempel vill att ditt fotohanteringsprogram ska starta när du ansluter en digitalkamera. Du kan också stänga av det här, så att inget händer när något ansluts.</p>
<p class="p">För att avgöra vilket program som ska startas när du ansluter olika enheter:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ikonen längst till höger i <span class="gui">menyraden</span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="guiseq"><span class="gui">Detaljer</span> ▸ <span class="gui">Flyttbar media</span></span>.</p></li>
<li class="steps">
<p class="p">Hitta din enhet eller mediatyp och välj sedan ett program eller en åtgärd för den mediatypen. Se nedan för en beskrivning av de olika typerna av enheter och media.</p>
<p class="p">Istället för att starta ett program kan du också ställa in att enheten ska visas i filhanteraren. När det händer kommer du tillfrågas om en åtgärd, annars händer inget automatiskt.</p>
</li>
<li class="steps"><p class="p">Alternativet <span class="gui">Mjukvara</span> skiljer sig lite från de övriga - om datorn känner av att det finns mjukvara på en skiva som du matar in kan den försöka köra mjukvaran automatiskt om du vill. Detta är bra om du har ett program som är installerat på en CD och du vill starta det när skivan matas in (exempelvis ett bildspel).</p></li>
<li class="steps"><p class="p">Om du inte ser enheten eller mediatypen du vill ändra i listan (som Blu-ray-skivor eller e-bokläsare), klicka på <span class="gui">Övrig media</span> för att se en mer detaljerad lista över enheter. Välj typen av enhet eller media från den utfällbara listan <span class="gui">Typ</span> och program eller åtgärd från listan <span class="gui">Åtgärd</span>.</p></li>
</ol></div></div></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du inte vill att något program öppnas automatiskt, oavsett vad du ansluter, välj <span class="gui">Fråga aldrig eller starta aldrig program vid inmatning av media</span> längst ner i fönstret Flyttbara enheter.</p></div></div></div></div>
</div>
<div id="files-types-of-devices" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Typer av enheter och media</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Musikskivor</dt>
<dd class="terms"><p class="p">Välj det musikprogram eller ljudkopieringsprogram du tycker bäst om för att hantera cd-skivor. Om du använder musik-dvd (DVD-A), välj hur du vill öppna dem under <span class="gui">Övrig media</span>. Om du öppnar en musikskiva med filhanteraren kommer spåren visas som WAV-filer som du kan spela upp i valfritt musikprogram.</p></dd>
<dt class="terms">Videoskivor</dt>
<dd class="terms"><p class="p">Välj det filmprogram du tycker bäst om för att hantera dvd-filmer. Använd knappen <span class="gui">Övrig media</span> för att ange ett program för Blu-ray, HD DVD, video-cd (VCD), och super video-cd (SVCD). Om dvd-skivor eller andra videoskivor inte fungerar korrekt när du matar in dem, se <span class="link"><a href="video-dvd.html" title="Why won't DVDs play?">Why won't DVDs play?</a></span>.</p></dd>
<dt class="terms">Tomma skivor</dt>
<dd class="terms"><p class="p">Använd knappen <span class="gui">Övrig media</span> för att välja ett skivbrännarprogram för tomma CD-skivor, DVD-skivor, Blu-ray-skivor, och HD DVD-skivor.</p></dd>
<dt class="terms">Kameror och foton</dt>
<dd class="terms">
<p class="p">Använd den utfällbara menyn <span class="gui">Foton</span> för att välja ett fotohanteringsprogram som ska köras när du ansluter din digitalkamera, eller när du matar in ett mediakort från en kamera, som CF-, SD-, MMC-, eller MS-kort. Du kan också utan problem bläddra bland dina foton i filhanteraren.</p>
<p class="p">Under <span class="gui">Övrig media</span> kan du välja ett program för att öppna Kodaks bildskivor, som du kan få tillverkade i en butik. Dessa är vanliga CD-skivor med JPEG-bilder i en mapp med namnet <span class="file">PICTURES</span>.</p>
</dd>
<dt class="terms">Musikspelare</dt>
<dd class="terms"><p class="p">Välj ett program för att hantera musikbiblioteket på din bärbara musikspelare, eller hantera filerna själv med filhanteraren.</p></dd>
<dt class="terms">E-bokläsare</dt>
<dd class="terms"><p class="p">Använd knappen <span class="gui">Övrig media</span> för att välja ett program för att hantera böckerna på din e-bokläsare, eller hantera filerna själv med filhanteraren.</p></dd>
<dt class="terms">Programvara</dt>
<dd class="terms">
<p class="p">Vissa skivor och flyttbar media innehåller programvara som är tänkt att köras automatiskt när mediet matas in. Använd alternativet <span class="gui">Programvara</span> för att styra vad som händer när media med självstartande program matas in. Du kommer alltid tillfrågas om bekräftelse innan program körs.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">Kör aldrig programvara från media du inte litar på.</p></div></div></div></div>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="files.html#removable" title="Flyttbara enheter och externa diskar">Flyttbara enheter och externa diskar</a></li>
<li class="links "><a href="media.html#photos" title="Foton och digitalkameror">Foton</a></li>
<li class="links "><a href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a></li>
<li class="links "><a href="media.html#videos" title="Videor och videokameror">Videor</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
