<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Kontrollera hur mycket diskutrymme som finns kvar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="disk.html" title="Hårddiskar &amp; lagring">Hårddiskar &amp; lagring</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Kontrollera hur mycket diskutrymme som finns kvar</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Du kan kontrollera hur mycket diskutrymme som finns kvar med <span class="app">Diskanvändningsanalys</span> eller <span class="app">Systemövervakaren</span>.</p></div>
<div id="disk-usage-analyzer" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kontrollera med Diskanvändningsanalys</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att kontrollera ledigt diskutrymme och diskkapacitet med <span class="app">Diskanvändningsanalys</span>:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Öppna programmet <span class="app">Diskanvändningsanalysator</span> från <span class="gui">Dash</span>. Fönstret kommer visa <span class="gui">Total filsystemskapacitet</span> och <span class="gui">Total filsystemsanvändning</span>.</p></li>
<li class="list"><p class="p">Klicka på en av knapparna på verktygsraden och välj <span class="gui">Skanna Hem</span>, <span class="gui">Skanna filsystem</span>, <span class="gui">Skanna mapp</span>, eller <span class="gui">Skanna fjärrmapp</span>.</p></li>
</ul></div></div></div>
<p class="p">Informationen sorteras efter <span class="gui">Mapp</span>, <span class="gui">Användning</span>, <span class="gui">Storlek</span> och <span class="gui">Innehåll</span>. Se fler detaljer i <span class="link"><a href="https://help.gnome.org/users/baobab/stable/" title="https://help.gnome.org/users/baobab/stable/"><span class="app">Diskanvändningsanalys</span></a></span>.</p>
</div></div>
</div></div>
<div id="system-monitor" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kontrollera med Systemövervakaren</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att kontrollera ledigt diskutrymme och diskkapacitet med <span class="app">Systemövervakaren</span>:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna programmet <span class="app">Systemövervakaren</span> från <span class="gui">Dash</span>.</p></li>
<li class="steps"><p class="p">Välj fliken <span class="gui">Filsystem</span> för att se systemets partitioner och diskanvändning. Informationen sorteras efter <span class="gui">Totalt</span>, <span class="gui">Ledigt</span>, <span class="gui">Tillgängligt</span> och <span class="gui">Använt</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="disk-full" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Vad gör jag om disken är full?</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Om disken är full bör du:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Radera filer som inte behövs eller som du inte kommer använda mer.</p></li>
<li class="list"><p class="p">Gär en <span class="link"><a href="backup-why.html" title="Säkerhetskopiera dina viktiga filer">säkerhetskopia</a></span> av viktiga filer som du inte behöver för en tid framöver och ta bort dem från hårddisken.</p></li>
</ul></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="disk.html" title="Hårddiskar &amp; lagring">Hårddiskar &amp; lagring</a><span class="desc"> — <span class="link"><a href="disk-capacity.html" title="Kontrollera hur mycket diskutrymme som finns kvar">Diskutrymme</a></span>, <span class="link"><a href="disk-benchmark.html" title="Testa din hårddisks prestanda">prestanda</a></span>, <span class="link"><a href="disk-check.html" title="Kontrollera din hårddisk för problem">problem</a></span>, <span class="link"><a href="disk-partitions.html" title="Hantera volymer och partitioner">volymer och partitioner</a></span>...</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
