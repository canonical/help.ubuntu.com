<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Inställningar för användare och system</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Inställningar för användare och system</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-grid ">
<div class="links-grid-link"><a href="user-accounts.html" title="Användarkonton">Användarkonton</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="user-add.html" title="Add a new user account">Add user</a></span> or
      <span class="link"><a href="shell-guest-session.html" title="Launch a restricted guest session">guest user</a></span>,
      <span class="link"><a href="user-changepassword.html" title="Välj ditt lösenord">change password</a></span>,
      <span class="link"><a href="user-admin-change.html" title="Change who has administrative privileges">administrators</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="clock.html" title="Datum &amp; tid">Datum &amp; tid</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="clock-set.html" title="Ändra tid och datum">Ange datum och tid</a></span>, <span class="link"><a href="clock-timezone.html" title="Visa andra tidszoner">tidszon</a></span>, <span class="link"><a href="clock-calendar.html" title="Kalendermöten">kalender och möten</a></span>...</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="color.html" title="Hantera färginställningar">Hantera färginställningar</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="color-whyimportant.html" title="Varför är färghantering viktigt?">Varför är det här viktigt</a></span>, <span class="link"><a href="color.html#profiles" title="Färgprofiler">Färgprofiler</a></span>, <span class="link"><a href="color.html#calibration" title="Kalibrering">Hur man kalibrerar en enhet</a></span>...</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="media.html#sound" title="Grundinställningar ljud">Ljud</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="sound-volume.html" title="Change the sound volume">Volym</a></span>, <span class="link"><a href="sound-usespeakers.html" title="Use different speakers or headphones">högtalare och hörlurar</a></span>, <span class="link"><a href="sound-usemic.html" title="Använd en annan mikrofon">mikrofoner</a></span>...</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="mouse.html" title="Mus">Mus</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="mouse-lefthanded.html" title="Använd din mus som vänsterhänt">Vänsterhänt</a></span>, <span class="link"><a href="mouse-sensitivity.html" title="Justera hastigheten för musen och styrplattan">hastighet och känslighet</a></span>, <span class="link"><a href="mouse-touchpad-click.html" title="Klicka, dra, eller rulla med styrplattan">styrplatteklick och rullning</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="accounts.html" title="Nätkonton">Nätkonton</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="accounts-add.html" title="Lägg till ett konto">Lägg till kontakter, </a></span> <span class="link"><a href="accounts-remove.html" title="Ta bort ett konto">Ta bort konton, </a></span> <span class="link"><a href="accounts-disable-service.html" title="Avaktivera kontotjänster">Avaktivera tjänster</a></span></span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="power.html" title="På/av &amp; batteri">På/av &amp; batteri</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="power-suspend.html" title="What happens when I suspend my computer?">Suspend</a></span>,
      <span class="link"><a href="power-batterylife.html" title="Use less power and improve battery life">energy savings</a></span>,
      <span class="link"><a href="shell-exit.html#shutdown" title="Power off or restart">power off</a></span>,
      <span class="link"><a href="power-whydim.html" title="Why does my screen go dim after a while?">screen dimming</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="prefs-language.html" title="Region &amp; språk">Region &amp; språk</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="prefs-language-install.html" title="Install languages">Install languages</a></span>,
      <span class="link"><a href="session-language.html" title="Change which language you use">change language</a></span>,
      <span class="link"><a href="session-formats.html" title="Change date and measurement formats">region and formats</a></span>,
      <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">input sources</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">Indatakällor</a></span>, <span class="link"><a href="keyboard-cursor-blink.html" title="Gör att tangentbordsmarkören blinkar">blinkande markör</a></span>, <span class="link"><a href="windows-key.html" title='Vad är "Superknappen"?'>supertangent</a></span>, <span class="link"><a href="a11y.html#mobility" title="Rörelsehinder">tangentbordsåtkomst</a></span>...</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="prefs-display.html" title="Visning och skärm">Visning och skärm</a></div>
<div class="desc"><span class="desc">
      <span class="link"><a href="look-background.html" title="Byt skrivbordsbakgrund">Background</a></span>,
      <span class="link"><a href="look-resolution.html" title="Ändra storlek och rotation för skärmen">size and rotation</a></span>,
      <span class="link"><a href="display-dimscreen.html" title="Ställ in skärmens ljusstyrka">brightness</a></span>…
    </span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="wacom.html" title="Wacom Graphics Tablet">Wacom Graphics Tablet</a></div>
<div class="desc"><span class="desc">Adjust the settings of your Wacom tablet.</span></div>
</div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
