<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Tidssynkronisering med NTP</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="networking.html" title="Nätverk">Nätverk</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="dhcp.html" title="Dynamic Host Configuration Protocol (DHCP)">Föregående</a><a class="nextlinks-next" href="dm-multipath-chapter.html" title="DM-Multipath">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Tidssynkronisering med NTP</h1></div>
<div class="region">
<div class="contents">
<p class="para">NTP är ett TCP/IP protokoll för synkronisering av tid över ett nätverk. I grund och botten är det en klient som frågar en server efter nuvarande tid och använder det för att ställa in sin egen klocka.</p>
<p class="para">
Behind this simple description, there is a lot of complexity - there are tiers of NTP servers, with the tier one NTP servers connected to atomic clocks, and tier two and three servers spreading the load of actually handling requests across the Internet. Also the client software is a lot more complex than you might think - it has to factor out communication delays, and adjust the time in a way that does not upset all the other processes that run on the server. But luckily all that complexity is hidden from you! 
</p>
<p class="para">
Ubuntu uses ntpdate and ntpd. 
</p>
</div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="NTP.html#ntpdate" title="ntpdate">ntpdate</a></li>
<li class="links"><a class="xref" href="NTP.html#ntpd" title="ntpd">ntpd</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-installation" title="Installation">Installation</a></li>
<li class="links"><a class="xref" href="NTP.html#timeservers" title="Konfiguration">Konfiguration</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-status" title="View status">View status</a></li>
<li class="links"><a class="xref" href="NTP.html#ntp-references" title="Referenser">Referenser</a></li>
</ul></div>
<div class="sect2 sect" id="ntpdate"><div class="inner">
<div class="hgroup"><h2 class="title">ntpdate</h2></div>
<div class="region"><div class="contents">
<p class="para">
Ubuntu comes with ntpdate as standard, and will run it once at boot time to set up your time according to Ubuntu's NTP server.
</p>
<div class="code"><pre class="contents ">ntpdate -s ntp.ubuntu.com
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="ntpd"><div class="inner">
<div class="hgroup"><h2 class="title">ntpd</h2></div>
<div class="region"><div class="contents"><p class="para">
   The ntp daemon ntpd calculates the drift of your system clock and continuously adjusts it, so there are no large corrections that could 
   lead to inconsistent logs for instance. The cost is a little processing power and memory, but for a modern server this is negligible. 
   </p></div></div>
</div></div>
<div class="sect2 sect" id="ntp-installation"><div class="inner">
<div class="hgroup"><h2 class="title">Installation</h2></div>
<div class="region"><div class="contents">
<p class="para">
   To install ntpd, from a terminal prompt enter: 
   </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt-get install ntp</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="timeservers"><div class="inner">
<div class="hgroup"><h2 class="title">Konfiguration</h2></div>
<div class="region"><div class="contents">
<p class="para">
  Edit <span class="file filename">/etc/ntp.conf</span> to add/remove server lines.
  By default these servers are configured:
  </p>
<div class="code"><pre class="contents "># Use servers from the NTP Pool Project. Approved by Ubuntu Technical Board
# on 2011-02-08 (LP: #104525). See http://www.pool.ntp.org/join.html for
# more information.
server 0.ubuntu.pool.ntp.org
server 1.ubuntu.pool.ntp.org
server 2.ubuntu.pool.ntp.org
server 3.ubuntu.pool.ntp.org
</pre></div>
<p class="para">
	  After changing the config file you have to reload the
          <span class="app application">ntpd</span>:
	  </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo service ntp reload</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="ntp-status"><div class="inner">
<div class="hgroup"><h2 class="title">View status</h2></div>
<div class="region"><div class="contents">
<p class="para">
  Use ntpq to see more info: 
  </p>
<div class="screen"><pre class="contents "><span class="cmd command"># sudo ntpq -p</span>
<span class="output computeroutput">     remote           refid      st t when poll reach   delay   offset  jitter
==============================================================================
+stratum2-2.NTP. 129.70.130.70    2 u    5   64  377   68.461  -44.274 110.334
+ntp2.m-online.n 212.18.1.106     2 u    5   64  377   54.629  -27.318  78.882
*145.253.66.170  .DCFa.           1 u   10   64  377   83.607  -30.159  68.343
+stratum2-3.NTP. 129.70.130.70    2 u    5   64  357   68.795  -68.168 104.612
+europium.canoni 193.79.237.14    2 u   63   64  337   81.534  -67.968  92.792</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="ntp-references"><div class="inner">
<div class="hgroup"><h2 class="title">Referenser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
  	    <p class="para">
          See the <a href="https://help.ubuntu.com/community/UbuntuTime" class="ulink" title="https://help.ubuntu.com/community/UbuntuTime">Ubuntu Time</a> wiki page for more information.
        </p>
      </li>
<li class="list itemizedlist">
  	    <p class="para">
          <a href="http://www.ntp.org/" class="ulink" title="http://www.ntp.org/">ntp.org, home of the Network Time Protocol project</a>
        </p>
      </li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="dhcp.html" title="Dynamic Host Configuration Protocol (DHCP)">Föregående</a><a class="nextlinks-next" href="dm-multipath-chapter.html" title="DM-Multipath">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
