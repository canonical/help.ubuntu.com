<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Handbok för Ubuntu-skrivbordet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" class="media media-inline" alt="Ubuntus logotyp"></span></span> Handbok för Ubuntu-skrivbordet</span></h1></div>
<div class="title" style="margin-bottom: 1.5em"><span>Ubuntu 18.04</span></div><div class="region"><div class="contents">
<div class="links topiclinks"><div class="inner"><div class="region"><div class="linkdiv "><a class="linkdiv" href="getting-started.html.sv" title="Komma igång"><span class="title">Börja med GNOME</span><span class="linkdiv-dash"> — </span><span class="desc">Är GNOME nytt för dig? Lär dig hur du använder det.</span></a></div></div></div></div>
<div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="shell-introduction.html.sv" title="Introduktion till GNOME"><span class="title">Introduktion till GNOME</span><span class="linkdiv-dash"> — </span><span class="desc">En visuell introduktion till ditt skrivbord, systemraden, och översiktsvyn <span class="gui">Aktiviteter</span>.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-exit.html.sv" title="Logga ut, stäng av eller växla användare"><span class="title">Logga ut, stäng av eller växla användare</span><span class="linkdiv-dash"> — </span><span class="desc">Lär dig hur du lämnar ditt användarkonto genom att logga ut, växla användare, och så vidare.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-apps-open.html.sv" title="Starta program"><span class="title">Starta program</span><span class="linkdiv-dash"> — </span><span class="desc">Starta program från översiktsvyn <span class="gui">Aktiviteter</span>.</span></a></div>
</div></div></div>
<div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-grid ">
<div class="links-grid-link"><a href="shell-overview.html.sv" title="Ditt skrivbord">Ditt skrivbord</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="clock-calendar.html.sv" title="Kalendermöten">Kalender</a></span>, <span class="link"><a href="shell-notifications.html.sv" title="Aviseringar och meddelandefältet">aviseringar</a></span>, <span class="link"><a href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar">tangentbordsgenvägar</a></span>, <span class="link"><a href="shell-windows.html.sv" title="Fönster och arbetsytor">fönster och arbetsytor</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlöst</a></span>, <span class="link"><a href="net-wired.html.sv" title="Trådbundna nätverk">trådbundet</a></span>, <span class="link"><a href="net-problem.html.sv" title="Nätverksproblem">anslutningsproblem</a></span>, <span class="link"><a href="net-browser.html.sv" title="Webbläsare">webbsurfning</a></span>, <span class="link"><a href="net-email.html.sv" title="E-post &amp; e-postprogramvara">e-postkonton</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="media.html.sv" title="Ljud, video och bilder">Ljud, video och bilder</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="media.html.sv#photos" title="Foton och digitalkameror">Digitalkameror</a></span>, <span class="link"><a href="media.html.sv#music" title="Musik och bärbara ljudspelare">iPod-enheter</a></span>, <span class="link"><a href="media.html.sv#photos" title="Foton och digitalkameror">redigera foton</a></span>, <span class="link"><a href="media.html.sv#videos" title="Videor och videokameror">spela upp videor</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="files.html.sv" title="Filer, mappar och sökning">Filer, mappar och sökning</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="files-search.html.sv" title="Sök efter filer">Sökning</a></span>, <span class="link"><a href="files-delete.html.sv" title="Ta bort filer och mappar">ta bort filer</a></span>, <span class="link"><a href="files.html.sv#backup" title="Säkerhetskopiering">säkerhetskopiering</a></span>, <span class="link"><a href="files.html.sv#removable" title="Flyttbara enheter och externa diskar">flyttbara enheter</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="addremove.html.sv" title="Installera &amp; ta bort mjukvara">Installera &amp; ta bort mjukvara</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="addremove-install.html.sv" title="Installera fler program">Installera program</a></span>, <span class="link"><a href="addremove-remove.html.sv" title="Ta bort ett program">ta bort program</a></span>, <span class="link"><a href="addremove-sources.html.sv" title="Lägg till fler programförråd">lägg till förråd</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="keyboard.html.sv" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html.sv" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html.sv" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html.sv" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html.sv" title="Användarkonton">användarkonton</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="hardware.html.sv" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="hardware.html.sv#problems" title="Vanliga problem">Hårdvaruproblem</a></span>, <span class="link"><a href="printing.html.sv" title="Utskrifter">skrivare</a></span>, <span class="link"><a href="power.html.sv" title="Ström och batteri">ströminställningar</a></span>, <span class="link"><a href="color.html.sv" title="Färghantering">färghantering</a></span>, <span class="link"><a href="bluetooth.html.sv" title="Bluetooth">Bluetooth</a></span>, <span class="link"><a href="disk.html.sv" title="Diskar och lagring">diskar</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="a11y.html.sv" title="Hjälpmedel">Hjälpmedel</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="a11y.html.sv#vision" title="Synnedsättningar">Se</a></span>, <span class="link"><a href="a11y.html.sv#sound" title="Hörselnedsättningar">höra</a></span>, <span class="link"><a href="a11y.html.sv#mobility" title="Rörelsehinder">mobilitet</a></span>, <span class="link"><a href="a11y-braille.html.sv" title="Läs skärmen med punktskrift">punktskrift</a></span>, <span class="link"><a href="a11y-mag.html.sv" title="Förstora en del av skärmen">skärmförstorare</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="tips.html.sv" title="Tips och tricks">Tips och tricks</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="tips-specialchars.html.sv" title="Mata in speciella tecken">Specialtecken</a></span>, <span class="link"><a href="mouse-middleclick.html.sv" title="Mittenklick">genvägar för mittenklick</a></span>…</span></div>
</div>
<div class="links-grid ">
<div class="links-grid-link"><a href="more-help.html.sv" title="Få mer hjälp">Få mer hjälp</a></div>
<div class="desc"><span class="desc"><span class="link"><a href="about-this-guide.html.sv" title="Om denna handbok">Användningstips</a></span>, <span class="link"><a href="get-involved.html.sv" title="Medverka till att förbättra den här handboken">hjälp till att förbättra handboken</a></span>…</span></div>
</div>
</div></div></div>
</div></div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
