<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Hitta program, filer, musik med mera med Snabbstartspanelen</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Hitta program, filer, musik med mera med Snabbstartspanelen</span></h1></div>
<div class="region">
<div class="contents">
<div class="media media-image floatend"><div class="inner"><img src="figures/unity-dash-sample.png" class="media media-block" alt="Unity Sök"></div></div>
<p class="p"><span class="gui">Snabbstartspanelen</span> låter dig söka efter program, filer, musik, och videor, och visar dig objekt som du har använt nyligen. Om du någonsin arbetat med ett kalkylark eller redigerat en bild och glömt var de har sparats kommer du helt säkert uppskatta den här funktionen i Snabbstartspanelen.</p>
<p class="p">För att börja använda <span class="gui">Snabbstartspanelen</span>, klicka på den övre ikonen i <span class="link"><a href="unity-launcher-intro.html" title="Använda programstartaren">Startaren</a></span>. Den här ikonen visar Ubuntus logo. För snabbare åtkomst kan du också trycka på <span class="key"><a href="windows-key.html" title='Vad är "Superknappen"?'><kbd>Supertangenten</kbd></a></span>.</p>
<p class="p">För att dölja <span class="gui">Snabbstartspanelen</span>, klicka på den övre ikonen igen, eller tryck <span class="key"><kbd>Super</kbd></span> eller <span class="key"><kbd>Esc</kbd></span>.</p>
</div>
<div id="dash-home" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Sök efter allt från Snabbstartspanelens hem</span></h2></div>
<div class="region">
<div class="contents">
<p class="p">Det första du ser när du öppnar Snabbstartspanelen är dess hemsida. Utan att skriva eller klicka på något kommer Snabbstartspanelens Hem visa dig program och filer som du använt nyligen.</p>
<p class="p">Bara en rad med resultat kommer visas för varje typ. Om det finns fler resultat kan du klicka på <span class="gui">Se fler resultat</span> för att se dem.</p>
<p class="p">För att söka, börja bara skriva så kommer möjliga sökträffar dyka upp automatiskt från de olika installerade linserna.</p>
<p class="p">Klicka på ett resultat för att öppna det, eller tryck <span class="key"><kbd>Retur</kbd></span> för att öppna det första objektet i listan.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="unity-shopping.html" title="Varför finns det shoppinglänkar i Dash?">Varför finns det shoppinglänkar i Dash?</a><span class="desc"> — Online-resultat gör Snabbstartspanelen mer användbar, och hjälper till att finansiera Ubuntus utveckling.</span>
</li>
<li class="links ">
<a href="shell-apps-favorites.html" title="Ändra vilka program som visas i Startaren">Ändra vilka program som visas i Startaren</a><span class="desc"> — Lägg till, flytta, eller ta bort ofta använda programikoner på Startaren.</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="dash-lenses" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Vyer</span></h2></div>
<div class="region">
<div class="contents">
<p class="p">Linser låter dig fokusera Snabbstartspanelens resultat, och exkludera resultat från andra linser.</p>
<p class="p">Du kan se de tillgängliga linserna i <span class="gui">linsraden</span>, den mörkare remsan längst ner i Snabbstartspanelen.</p>
<p class="p">För att växla till en annan lins, klicka på den relevanta ikonen eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span>.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul>
<li class="links ">
<a href="unity-dash-files.html" title="Filvy">Filvy</a><span class="desc"> — Hitta filer, mappar, och nedladdningar.</span>
</li>
<li class="links ">
<a href="unity-dash-photos.html" title="Fotolinsen">Fotolinsen</a><span class="desc"> — Visa bilder från din dator eller dina sociala medier.</span>
</li>
<li class="links ">
<a href="unity-dash-music.html" title="Musiklins">Musiklins</a><span class="desc"> — Hitta och spela musik från din dator eller från internet.</span>
</li>
<li class="links ">
<a href="unity-dash-apps.html" title="Programlins">Programlins</a><span class="desc"> — Kör, installera, eller avinstallera program.</span>
</li>
<li class="links ">
<a href="unity-dash-video.html" title="Videolins">Videolins</a><span class="desc"> — Hitta och spela upp videor från din dator eller internet.</span>
</li>
<li class="links ">
<a href="unity-dash-friends.html" title="Vänner">Vänner</a><span class="desc"> — Bläddra bland meddelanden från dina konton hos sociala medier.</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="dash-filters" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Filter</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Filter låter dig begränsa din sökning ännu mer.</p>
<p class="p">Klicka på <span class="gui">Filtrera resultat</span> för att välja filter. Du kan behöva klicka på en filterrubrik, som <span class="gui">Källor</span> för att se möjliga alternativ.</p>
</div></div>
</div></div>
<div id="dash-previews" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Förhandsvisningar</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Om du högerklickar på ett sökresultat kommer en <span class="gui">förhandsgranskning</span> öppnas med mer information om sökresultatet.</p>
<p class="p">För att stänga förhandsgranskningen, klicka på en tom yta eller tryck <span class="key"><kbd>Esc</kbd></span>.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
