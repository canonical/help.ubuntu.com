<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Byt namn på en fil eller mapp</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#common-file-tasks" title="Vanliga åtgärder">Vanliga åtgärder</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Byt namn på en fil eller mapp</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Som med andra filhanterare kan du använda <span class="app">Filer</span> för att byta namn på en fil eller mapp.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">För att byta namn på en fil eller mapp:</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Högerklicka på objektet och välj <span class="gui">Byt namn</span> eller markera filen och tryck på <span class="key"><kbd>F2</kbd></span>.</p></li>
<li class="steps"><p class="p">Ange det nya namnet och tryck på <span class="key"><kbd>Retur</kbd></span> eller klicka på <span class="gui">Byt namn</span>.</p></li>
</ol></div>
</div></div>
<p class="p">Du kan också byta namn på en fil från fönstret<span class="link"><a href="nautilus-file-properties-basic.html.sv" title="Filegenskaper">egenskaper</a></span>.</p>
<p class="p">När du byter namn på en fil kommer bara första delen av namnet på filen att markeras, inte filändelsen (delen efter sista <span class="file">.</span>). Filändelsen betecknar vanligtvis vilken typ av fil det är (till exempel är <span class="file">file.pdf</span> ett PDF-dokument) och du vill vanligtvis inte ändra den. Om du behöver ändra filändelsen också så välj hela filnamnet och ändra det.</p>
<div class="note note-tip" title="Tips">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m12 2c-3.8541 0-7 3.1459-7 7 0 1.823 0.4945 3.139 1.1641 4.133 0.6695 0.994 1.4328 1.671 2.039 2.471 0.0882 0.116 0.1749 0.656 0.2071 1.32 0.016 0.332 0.0133 0.68 0.1894 1.119 0.0881 0.22 0.2439 0.478 0.5059 0.672 0.2619 0.194 0.6028 0.285 0.8945 0.285h4c0.583 0 1.204-0.478 1.402-0.908 0.199-0.43 0.217-0.793 0.244-1.137 0.056-0.688 0.138-1.319 0.211-1.441 0.549-0.916 1.304-2.009 1.94-3.114 0.636-1.104 1.203-2.199 1.203-3.4 0-3.8541-3.146-7-7-7zm0 2c2.773 0 5 2.2267 5 5 0 0.456-0.359 1.401-0.936 2.402-0.111 0.195-0.246 0.399-0.369 0.598h-7.8825c-0.4871-0.728-0.8125-1.519-0.8125-3 0-2.7733 2.2267-5 5-5z" style="block-progression:tb;color-rendering:auto;color:#000000;image-rendering:auto;isolation:auto;mix-blend-mode:normal;shape-rendering:auto;solid-color:#000000;text-decoration-color:#000000;text-decoration-line:none;text-decoration-style:solid;text-indent:0;text-transform:none;white-space:normal"></path>
 <path class="yelp-svg-fill" d="m9 20a0.5 0.5 0 0 0-0.5 0.5 0.5 0.5 0 0 0 0.5 0.5h6a0.5 0.5 0 0 0 0.5-0.5 0.5 0.5 0 0 0-0.5-0.5h-6zm0 2a0.5 0.5 0 0 0-0.5 0.5 0.5 0.5 0 0 0 0.5 0.5h6a0.5 0.5 0 0 0 0.5-0.5 0.5 0.5 0 0 0-0.5-0.5h-6z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Om du bytt namn på fel fil eller gav filen fel namn kan du ångra namnbytet. För att ångra åtgärden tryck omedelbart på menyknappen i verktygsfältet och välj <span class="gui">Ångra namnbyte</span>, eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Z</kbd></span></span> för att återställa det gamla namnet.</p></div></div></div>
</div>
</div>
<section id="valid-chars"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Giltiga tecken för filnamn</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Du kan använda vilket tecken som helst i filnamn förutom tecknet <span class="file">/</span> (snedstreck). Vissa enheter använder dock ett <span class="em">filsystem</span> som har fler restriktioner på filnamnen. Därför är det bäst att undvika följande tecken i dina filnamn: <span class="file">|</span>, <span class="file">\</span>, <span class="file">?</span>, <span class="file">*</span>, <span class="file">&lt;</span>, <span class="file">"</span>, <span class="file">:</span>, <span class="file">&gt;</span>, <span class="file">/</span>.</p>
<div class="note note-warning" title="Varning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m11.92 3.3047a1.3872 1.3872 0 0 0-1.129 0.6933l-8.6055 14.922a1.3872 1.3872 0 0 0 1.2012 2.08l17.226-8e-3a1.3872 1.3872 0 0 0 1.201-2.08l-8.619-14.916a1.3872 1.3872 0 0 0-1.136-0.6913 1.3872 1.3872 0 0 0-0.139 0zm0.08 4.6953a1 1 0 0 1 1 1v6a1 1 0 0 1-1 1 1 1 0 0 1-1-1v-6a1 1 0 0 1 1-1zm0 9a1 1 0 0 1 1 1 1 1 0 0 1-1 1 1 1 0 0 1-1-1 1 1 0 0 1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Om du namnger en fil med en <span class="file">.</span> som första tecken kommer filen att bli <span class="link"><a href="files-hidden.html.sv" title="Dölj en fil">dold</a></span> när du försöker visa den i filhanteraren.</p></div></div></div>
</div>
</div></div>
</div></section><section id="common-probs"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Vanliga problem</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Filnamnet används redan</dt>
<dd class="terms">
<p class="p">Du kan inte ha två filer eller mappar med samma namn i samma mapp. Om du försöker att byta namn på en fil till ett namn som redan existerar i mappen du arbetar i kommer filhanteraren inte att tillåta det.</p>
<p class="p">Fil- och mappnamn är skiftlägeskänsliga, så filnamnet <span class="file">File.txt</span> är inte detsamma som <span class="file">FILE.txt</span>. Att använda olika filnamn på detta sätt är tillåtet, men det är inte rekommenderat.</p>
</dd>
<dt class="terms">Filnamnet är för långt</dt>
<dd class="terms"><p class="p">På vissa filsystem kan filnamn inte har mer än 255 tecken. Denna 255-teckensbegränsning inkluderar både filnamnet och sökvägen till filen (till exempel <span class="file">/home/maria/Dokument/arbete/affärsförslag/…</span>), så du bör undvika långa fil- och mappnamn där det går.</p></dd>
<dt class="terms">Alternativet att byta namn är inaktiverat</dt>
<dd class="terms"><p class="p">Om <span class="gui">Byt namn</span> är inaktiverat har du inte rättighet att byta namn på filen. Du bör vara aktsam med att byta namn på sådana filer, eftersom namnbyte på vissa skyddade filer kan orsaka att systemet blir instabilt. Se <span class="link"><a href="nautilus-file-properties-permissions.html.sv" title="Ange filrättigheter">Ange filrättigheter</a></span> för vidare information.</p></dd>
</dl></div></div></div></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html.sv#common-file-tasks" title="Vanliga åtgärder">Vanliga åtgärder</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
