<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Samba och LDAP</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="network-authentication.html" title="Nätverksautentisering">Nätverksautentisering</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="openldap-server.html" title="OpenLDAP-server">Föregående</a><a class="nextlinks-next" href="kerberos.html" title="Kerberos">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Samba och LDAP</h1></div>
<div class="region">
<div class="contents"><p class="para">
	This section covers the integration of Samba with LDAP. The Samba server's role will be that of a "standalone" server and the LDAP
	directory will provide the authentication layer in addition to containing the user, group, and machine account information that Samba
	requires in order to function (in any of its 3 possible roles). The pre-requisite is an OpenLDAP server configured with a directory
	that can accept authentication requests. See <a class="xref" href="openldap-server.html" title="OpenLDAP-server">OpenLDAP-server</a> for details on fulfilling this requirement. Once this
	section is completed, you will need to decide what specifically you want Samba to do for you and then configure it accordingly.
	</p></div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="samba-ldap.html#samba-ldap-installation" title="Software Installation">Software Installation</a></li>
<li class="links"><a class="xref" href="samba-ldap.html#samba-ldap-openldap-configuration" title="LDAP Configuration">LDAP Configuration</a></li>
<li class="links"><a class="xref" href="samba-ldap.html#samba-ldap-samba-configuration" title="Samba konfigurering">Samba konfigurering</a></li>
<li class="links"><a class="xref" href="samba-ldap.html#samba-ldap-resources" title="Resurser">Resurser</a></li>
</ul></div>
<div class="sect2 sect" id="samba-ldap-installation"><div class="inner">
<div class="hgroup"><h2 class="title">Software Installation</h2></div>
<div class="region"><div class="contents">
<p class="para">
	There are three packages needed when integrating Samba with LDAP: <span class="app application">samba</span>, <span class="app application">samba-doc</span>,
	and <span class="app application">smbldap-tools</span> packages.
	</p>
<p class="para">
	Strictly speaking, the <span class="app application">smbldap-tools</span> package isn't needed, but unless you have some other way to manage the various
	Samba entities (users, groups, computers) in an LDAP context then you should install it.  
	</p>
<p class="para">
	Install these packages now:
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt-get install samba samba-doc smbldap-tools</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="samba-ldap-openldap-configuration"><div class="inner">
<div class="hgroup"><h2 class="title">LDAP Configuration</h2></div>
<div class="region">
<div class="contents">
<p class="para">
	We will now configure the LDAP server so that it can accomodate Samba data. We will perform three tasks in this section:
	</p>
<div class="steps"><div class="inner"><ol class="steps">
<li class="steps">
		<p class="para">Import a schema</p>
		</li>
<li class="steps">
		<p class="para">Index some entries</p>
		</li>
<li class="steps">
		<p class="para">Add objects</p>
		</li>
</ol></div></div>
</div>
<div class="sect3 sect" id="samba-ldap-openldap-configuration-samba-schema"><div class="inner">
<div class="hgroup"><h3 class="title">Samba schema</h3></div>
<div class="region"><div class="contents">
<p class="para">
      	In order for OpenLDAP to be used as a backend for Samba, logically, the DIT will need to use attributes that can properly describe
	Samba data. Such attributes can be obtained by introducing a Samba LDAP schema. Let's do this now.
      	</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
		<p class="para">
		For more information on schemas and their installation see <a class="xref" href="openldap-server.html#openldap-configuration" title="Modifying the slapd Configuration Database">Modifying the slapd Configuration Database</a>.
		</p>
	</div></div></div></div>
<div class="steps"><div class="inner"><ol class="steps">
<li class="steps">
		<p class="para">
		The schema is found in the now-installed <span class="app application">samba-doc</span> package. It needs to be unzipped and copied to 
		the <span class="file filename">/etc/ldap/schema</span> directory:
		</p>
        
<div class="screen"><pre class="contents "><span class="cmd command">sudo cp /usr/share/doc/samba-doc/examples/LDAP/samba.schema.gz /etc/ldap/schema</span>
<span class="cmd command">sudo gzip -d /etc/ldap/schema/samba.schema.gz</span>
</pre></div>

	</li>
<li class="steps">
		<p class="para">                  
		Have the configuration file <span class="file filename">schema_convert.conf</span> that contains the following lines:
		</p>

<div class="code"><pre class="contents ">include /etc/ldap/schema/core.schema
include /etc/ldap/schema/collective.schema
include /etc/ldap/schema/corba.schema
include /etc/ldap/schema/cosine.schema
include /etc/ldap/schema/duaconf.schema
include /etc/ldap/schema/dyngroup.schema
include /etc/ldap/schema/inetorgperson.schema
include /etc/ldap/schema/java.schema
include /etc/ldap/schema/misc.schema
include /etc/ldap/schema/nis.schema
include /etc/ldap/schema/openldap.schema
include /etc/ldap/schema/ppolicy.schema
include /etc/ldap/schema/ldapns.schema
include /etc/ldap/schema/pmi.schema
include /etc/ldap/schema/samba.schema
</pre></div>

	</li>
<li class="steps">
                <p class="para">
                Have the directory <span class="file filename">ldif_output</span> hold output.
                </p> 
       	</li>
<li class="steps">
		<p class="para">
		Determine the index of the schema:
		</p>

<div class="screen"><pre class="contents "><span class="cmd command">slapcat -f schema_convert.conf -F ldif_output -n 0 | grep samba,cn=schema</span>
<span class="output computeroutput">
dn: cn={14}samba,cn=schema,cn=config
</span>
</pre></div>

	</li>
<li class="steps">
                <p class="para">
                Convert the schema to LDIF format:
                </p>

<div class="screen"><pre class="contents "><span class="cmd command">slapcat -f schema_convert.conf -F ldif_output -n0 -H \
ldap:///cn={14}samba,cn=schema,cn=config -l cn=samba.ldif</span>
</pre></div>

       	</li>
<li class="steps">
                <p class="para">
                Edit the generated <span class="file filename">cn=samba.ldif</span> file by removing index information to arrive at:
                </p> 

<div class="code"><pre class="contents ">dn: cn=samba,cn=schema,cn=config
...
cn: samba
</pre></div>
		
                <p class="para">
                Remove the bottom lines:
                </p> 

<div class="code"><pre class="contents ">structuralObjectClass: olcSchemaConfig
entryUUID: b53b75ca-083f-102d-9fff-2f64fd123c95
creatorsName: cn=config
createTimestamp: 20080827045234Z
entryCSN: 20080827045234.341425Z#000000#000#000000
modifiersName: cn=config
modifyTimestamp: 20080827045234Z
</pre></div>

		<p class="para">
		Your attribute values will vary.
		</p>
	</li>
<li class="steps">
                <p class="para">
                Add the new schema:
                </p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo ldapadd -Q -Y EXTERNAL -H ldapi:/// -f cn\=samba.ldif</span>
</pre></div>

                <p class="para">
                To query and view this new schema:
                </p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo ldapsearch -Q -LLL -Y EXTERNAL -H ldapi:/// -b cn=schema,cn=config 'cn=*samba*'</span>
</pre></div>

	</li>
</ol></div></div>
</div></div>
</div></div>
<div class="sect3 sect" id="samba-ldap-openldap-configuration-samba-indices"><div class="inner">
<div class="hgroup"><h3 class="title">Samba indices</h3></div>
<div class="region"><div class="contents">
<p class="para">
	Now that slapd knows about the Samba attributes, we can set up some indices based on them. Indexing entries is a way to improve
	performance when a client performs a filtered search on the DIT.
	</p>
<p class="para">
	Create the file <span class="file filename">samba_indices.ldif</span> with the following contents:
	</p>
<div class="code"><pre class="contents ">dn: olcDatabase={1}hdb,cn=config
changetype: modify
add: olcDbIndex
olcDbIndex: uidNumber eq
olcDbIndex: gidNumber eq
olcDbIndex: loginShell eq
olcDbIndex: uid eq,pres,sub
olcDbIndex: memberUid eq,pres,sub
olcDbIndex: uniqueMember eq,pres
olcDbIndex: sambaSID eq
olcDbIndex: sambaPrimaryGroupSID eq
olcDbIndex: sambaGroupType eq
olcDbIndex: sambaSIDList eq
olcDbIndex: sambaDomainName eq
olcDbIndex: default sub
</pre></div>
<p class="para">
	Using the <span class="app application">ldapmodify</span> utility load the new indices:
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo ldapmodify -Q -Y EXTERNAL -H ldapi:/// -f samba_indices.ldif</span>
</pre></div>
<p class="para">
	If all went well you should see the new indices using <span class="app application">ldapsearch</span>:
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo ldapsearch -Q -LLL -Y EXTERNAL -H \
ldapi:/// -b cn=config olcDatabase={1}hdb olcDbIndex</span>
</pre></div>
</div></div>
</div></div>
<div class="sect3 sect" id="samba-ldap-openldap-configuration-populating"><div class="inner">
<div class="hgroup"><h3 class="title">Adding Samba LDAP objects</h3></div>
<div class="region"><div class="contents">
<p class="para">
	Next, configure the <span class="app application">smbldap-tools</span> package to match your environment.  The package 
	is supposed to come with a configuration helper script (smbldap-config.pl, formerly configure.pl) that will ask questions
	about the needed options but there is a <a href="https://bugs.launchpad.net/serverguide/+bug/997172" class="ulink" title="https://bugs.launchpad.net/serverguide/+bug/997172">bug</a>
	whereby it is not installed (but found in the source code; 'apt-get source smbldap-tools').
	</p>
<p class="para">
	To manually configure the package, you need to create and edit the files <span class="file filename">/etc/smbldap-tools/smbldap.conf</span> and
	<span class="file filename">/etc/smbldap-tools/smbldap_bind.conf</span>.
	</p>
<p class="para">
	The <span class="app application">smbldap-populate</span> script will then add the LDAP objects required for Samba. It is a good idea to first
	make a backup of your DIT using <span class="app application">slapcat</span>:
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo slapcat -l backup.ldif</span>
</pre></div>
<p class="para">
	Once you have a backup proceed to populate your directory:
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo smbldap-populate</span>
</pre></div>
<p class="para">
	You can create a LDIF file containing the new Samba objects by executing <span class="cmd command">sudo smbldap-populate -e samba.ldif</span>.
	This allows you to look over the changes making sure everything is correct. If it is, rerun the script without the '-e'
	switch. Alternatively, you can take the LDIF file and import its data per usual.
	</p>
<p class="para">
	Your LDAP directory now has the necessary information to authenticate Samba users.
	</p>
</div></div>
</div></div>
</div>
</div></div>
<div class="sect2 sect" id="samba-ldap-samba-configuration"><div class="inner">
<div class="hgroup"><h2 class="title">Samba konfigurering</h2></div>
<div class="region"><div class="contents">
<p class="para">
	There are multiple ways to configure Samba. For details on some common configurations see <a class="xref" href="samba.html" title="Samba">Samba</a>.      
	To configure Samba to use LDAP, edit its configuration file <span class="file filename">/etc/samba/smb.conf</span> commenting out
	the default <span class="em emphasis">passdb backend</span> parameter and adding some ldap-related ones:
	</p>
<div class="code"><pre class="contents ">#   passdb backend = tdbsam

# LDAP Settings
   passdb backend = ldapsam:ldap://hostname
   ldap suffix = dc=example,dc=com
   ldap user suffix = ou=People
   ldap group suffix = ou=Groups
   ldap machine suffix = ou=Computers
   ldap idmap suffix = ou=Idmap
   ldap admin dn = cn=admin,dc=example,dc=com
   ldap ssl = start tls
   ldap passwd sync = yes
...
   add machine script = sudo /usr/sbin/smbldap-useradd -t 0 -w "%u"
</pre></div>
<p class="para">
	Change the values to match your environment.
	</p>
<p class="para">Starta om <span class="app application">samba</span> för att aktivera de nya inställningarna:</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo restart smbd</span>
<span class="cmd command">sudo restart nmbd</span>
</pre></div>
<p class="para">
	Now inform Samba about the rootDN user's password (the one set during the installation of the slapd package):
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo smbpasswd -w password</span>
</pre></div>
<p class="para">
	If you have existing LDAP users that you want to include in your new LDAP-backed Samba they will, of course, also need to be given
	some of the extra attributes. The <span class="app application">smbpasswd</span> utility can do this as well (your host will need to be
	able to see (enumerate) those users via NSS; install and configure either <span class="app application">libnss-ldapd</span> or
	<span class="app application">libnss-ldap</span>):
	</p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo smbpasswd -a användarnamn</span>
</pre></div>
<p class="para">
	You will prompted to enter a password. It will be considered as the new password for that user. Making it the same as before is reasonable.
	</p>
<p class="para">
	To manage user, group, and machine accounts use the utilities provided by the <span class="app application">smbldap-tools</span> package.
	Here are some examples:
	</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
		<p class="para">
		To add a new user:
		</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo smbldap-useradd -a -P användarnamn</span>
</pre></div>

		<p class="para">
		The <span class="em emphasis">-a</span> option adds the Samba attributes, and the <span class="em emphasis">-P</span> option calls the 
		<span class="app application">smbldap-passwd</span> utility after the user is created allowing you to enter a password for the user.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		To remove a user:
		</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo smbldap-userdel användarnamn</span>
</pre></div>

		<p class="para">
		In the above command, use the <span class="em emphasis">-r</span> option to remove the user's home directory.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		To add a group:
		</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo smbldap-groupadd -a gruppnamn</span>
</pre></div>

		<p class="para">
		As for <span class="app application">smbldap-useradd</span>, the <span class="em emphasis">-a</span> adds the Samba attributes.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		To make an existing user a member of a group:
		</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo smbldap-groupmod -m användarnamn gruppnamn</span>
</pre></div>

		<p class="para">
		The <span class="em emphasis">-m</span> option can add more than one user at a time by listing them in comma-separated format.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		To remove a user from a group:
		</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo smbldap-groupmod -x användarnamn gruppnamn</span>
</pre></div>

		</li>
<li class="list itemizedlist">
		<p class="para">
		To add a Samba machine account:
		</p>

<div class="screen"><pre class="contents "><span class="cmd command">sudo smbldap-useradd -t 0 -w användarnamn</span>
</pre></div>

		<p class="para">
		Replace <span class="em emphasis">username</span> with the name of the workstation.  The <span class="em emphasis">-t 0</span> option creates the machine account
		without a delay, while the <span class="em emphasis">-w</span> option specifies the user as a machine account.  Also, note the 
		<span class="em emphasis">add machine script</span> parameter in <span class="file filename">/etc/samba/smb.conf</span> was changed to use <span class="app application">smbldap-useradd</span>.
		</p>
		</li>
</ul></div>
<p class="para">
	There are utilities in the <span class="app application">smbldap-tools</span> package that were not covered here. Here is a complete list:
	</p>
<div class="code"><pre class="contents "><a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupadd.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupadd.8.html">smbldap-groupadd</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupdel.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupdel.8.html">smbldap-groupdel</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupmod.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupmod.8.html">smbldap-groupmod</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupshow.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-groupshow.8.html">smbldap-groupshow</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-passwd.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-passwd.8.html">smbldap-passwd</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-populate.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-populate.8.html">smbldap-populate</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-useradd.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-useradd.8.html">smbldap-useradd</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-userdel.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-userdel.8.html">smbldap-userdel</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-userinfo.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-userinfo.8.html">smbldap-userinfo</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-userlist.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-userlist.8.html">smbldap-userlist</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-usermod.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-usermod.8.html">smbldap-usermod</a>
<a href="http://manpages.ubuntu.com/manpages/en/man8/smbldap-usershow.8.html" class="ulink" title="http://manpages.ubuntu.com/manpages/en/man8/smbldap-usershow.8.html">smbldap-usershow</a>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="samba-ldap-resources"><div class="inner">
<div class="hgroup"><h2 class="title">Resurser</h2></div>
<div class="region"><div class="contents"><div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
		<p class="para">
		For more information on installing and configuring Samba see <a class="xref" href="samba.html" title="Samba">Samba</a> of this Ubuntu Server Guide.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		There are multiple places where LDAP and Samba is documented in the upstream
		<a href="http://samba.org/samba/docs/man/Samba-HOWTO-Collection/" class="ulink" title="http://samba.org/samba/docs/man/Samba-HOWTO-Collection/">Samba HOWTO Collection</a>.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		Regarding the above, see specifically the <a href="http://samba.org/samba/docs/man/Samba-HOWTO-Collection/passdb.html" class="ulink" title="http://samba.org/samba/docs/man/Samba-HOWTO-Collection/passdb.html">passdb section</a>.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		Although dated (2007), the <a href="http://download.gna.org/smbldap-tools/docs/samba-ldap-howto/" class="ulink" title="http://download.gna.org/smbldap-tools/docs/samba-ldap-howto/">Linux Samba-OpenLDAP HOWTO</a> contains valuable notes.
		</p>
		</li>
<li class="list itemizedlist">
		<p class="para">
		The main page of the <a href="https://help.ubuntu.com/community/Samba#samba-ldap" class="ulink" title="https://help.ubuntu.com/community/Samba#samba-ldap">Samba Ubuntu community documentation</a> has a plethora of links to
		articles that may prove useful.
		</p>
		</li>
</ul></div></div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="openldap-server.html" title="OpenLDAP-server">Föregående</a><a class="nextlinks-next" href="kerberos.html" title="Kerberos">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
