<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Starta program</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 19.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Starta program</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Flytta din musmarkör till <span class="gui">Aktiviteter</span> i övre vänstra hörnet på skärmen för att visa översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span>. Här kan du hitta alla dina program. Du kan också öppna översiktsvyn genom att trycka på tangenten <span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span>.</p>
<p class="p">Det finns flera sätt att öppna ett program när du väl är i översiktsvyn <span class="gui">Aktiviteter</span>:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Börja skriva namnet på ett program — sökningen börjar omedelbart. (Om detta inte händer klicka på sökraden i toppen på skärmen och börja skriv.) Om du inte känner till det exakta namnet på ett program, prova att skriva in en relaterad term. Klicka på programmets ikon för att starta det.</p></li>
<li class="list">
<p class="p">Vissa program har ikoner i <span class="em">snabbstartspanelen</span>, den vertikala raden av ikoner på vänster sida av översiktsvyn <span class="gui">Aktiviteter</span>. Klicka på en av dessa för att starta motsvarande program.</p>
<p class="p">Om du har program som du använder ofta kan du själv <span class="link"><a href="shell-apps-favorites.html.sv" title="Nåla fast dina favoritprogram i snabbstartspanelen">lägga till dem i snabbstartspanelen</a></span>.</p>
</li>
<li class="list"><p class="p">Klicka på rutnätsknappen längst ner i snabbstartspanelen. Du kommer att få se ofta använda program om vyn <span class="gui">Ofta använda</span> är aktiverad. Om du vill köra ett nytt program, tryck på knappen <span class="gui">Alla</span> längst ner för att visa alla programmen. Tryck på programmet för att starta det.</p></li>
<li class="list">
<p class="p">Du kan starta ett program i en separat <span class="link"><a href="shell-workspaces.html.sv" title="Vad är en arbetsyta, och hur hjälper den mig?">arbetsyta</a></span> genom att dra dess ikon från snabbstartspanelen och släppa den på en utav arbetsytorna på höger sida av skärmen. Programmet kommer att öppnas i den valda arbetsytan.</p>
<p class="p">Du kan starta ett program i en <span class="em">ny</span> arbetsyta genom dra dess ikon till den tomma arbetsytan längst ner i arbetsyteväxlaren, eller till det lilla mellanrummet mellan två arbetsytor.</p>
</li>
</ul></div></div></div>
<div class="note note-tip" title="Tips">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m12 2c-3.8541 0-7 3.1459-7 7 0 1.823 0.4945 3.139 1.1641 4.133 0.6695 0.994 1.4328 1.671 2.039 2.471 0.0882 0.116 0.1749 0.656 0.2071 1.32 0.016 0.332 0.0133 0.68 0.1894 1.119 0.0881 0.22 0.2439 0.478 0.5059 0.672 0.2619 0.194 0.6028 0.285 0.8945 0.285h4c0.583 0 1.204-0.478 1.402-0.908 0.199-0.43 0.217-0.793 0.244-1.137 0.056-0.688 0.138-1.319 0.211-1.441 0.549-0.916 1.304-2.009 1.94-3.114 0.636-1.104 1.203-2.199 1.203-3.4 0-3.8541-3.146-7-7-7zm0 2c2.773 0 5 2.2267 5 5 0 0.456-0.359 1.401-0.936 2.402-0.111 0.195-0.246 0.399-0.369 0.598h-7.8825c-0.4871-0.728-0.8125-1.519-0.8125-3 0-2.7733 2.2267-5 5-5z" style="block-progression:tb;color-rendering:auto;color:#000000;image-rendering:auto;isolation:auto;mix-blend-mode:normal;shape-rendering:auto;solid-color:#000000;text-decoration-color:#000000;text-decoration-line:none;text-decoration-style:solid;text-indent:0;text-transform:none;white-space:normal"></path>
 <path class="yelp-svg-fill" d="m9 20a0.5 0.5 0 0 0-0.5 0.5 0.5 0.5 0 0 0 0.5 0.5h6a0.5 0.5 0 0 0 0.5-0.5 0.5 0.5 0 0 0-0.5-0.5h-6zm0 2a0.5 0.5 0 0 0-0.5 0.5 0.5 0.5 0 0 0 0.5 0.5h6a0.5 0.5 0 0 0 0.5-0.5 0.5 0.5 0 0 0-0.5-0.5h-6z"></path>
</svg><div class="inner">
<div class="title title-note"><h2><span class="title">Kör ett kommando snabbt</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Ett annat sätt att start ett program är att trycka <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F2</kbd></span></span>, skriva in dess <span class="em">kommandonamn</span> och sedan trycka på <span class="key"><kbd>Retur</kbd></span>-tangenten.</p>
<p class="p">För att till exempel starta <span class="app">Rhythmbox</span>, tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F2</kbd></span></span> och skriv ”<span class="cmd">rhythmbox</span>” (utan citattecken). Namnet på programmet är kommandot som startar programmet.</p>
<p class="p">Använd piltangenterna för att snabbt komma åt tidigare körda kommandon.</p>
</div></div>
</div>
</div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="shell-overview.html.sv" title="Ditt skrivbord">Ditt skrivbord</a><span class="desc"> — <span class="link"><a href="clock-calendar.html.sv" title="Kalendermöten">Kalender</a></span>, <span class="link"><a href="shell-notifications.html.sv" title="Aviseringar och aviseringslistan">aviseringar</a></span>, <span class="link"><a href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar">tangentbordsgenvägar</a></span>, <span class="link"><a href="shell-windows.html.sv" title="Fönster och arbetsytor">fönster och arbetsytor</a></span>…</span>
</li>
<li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="gs-use-system-search.html.sv" title="Använd systemsökning">En handledning i att använda systemsökning</a></li>
<li class="links "><a href="gs-launch-applications.html.sv" title="Starta program">En handledning i att starta program</a></li>
<li class="links ">
<a href="shell-apps-favorites.html.sv" title="Nåla fast dina favoritprogram i snabbstartspanelen">Nåla fast dina favoritprogram i snabbstartspanelen</a><span class="desc"> — Lägg till (eller ta bort) ofta använda programikoner från snabbstartspanelen.</span>
</li>
</ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
