<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använda programstartaren</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Använda programstartaren</span></h1></div>
<div class="region">
<div class="contents">
<div class="media media-image floatstart"><div class="inner"><img src="figures/unity-launcher-apps.png" class="media media-block" alt="Launcher icons"></div></div>
<p class="p">The <span class="gui">Launcher</span> is one of the key components of the Unity desktop. When you log in
   to your desktop, it will appear along the left-hand side of the screen. The Launcher provides you
   with quick access to applications, workspaces, removable devices and the trash.</p>
<p class="p">If an application that you want to start using is present in the Launcher, you can click on that
   application's icon, and it will start up, ready for you to use.</p>
<p class="p">To learn more about the Launcher, explore any of the Launcher help topics below.</p>
</div>
<div id="launcher-using" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Use the Launcher</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="unity-launcher-menu.html" title="The Launcher Icon Menus"><span class="title">The Launcher Icon Menus</span><span class="linkdiv-dash"> — </span><span class="desc">Right clicking a Launcher Icon reveals a menu of actions.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-launcher-shapes.html" title="What do the different shapes and colors in Launcher icons mean?"><span class="title">What do the different shapes and colors in Launcher icons mean?</span><span class="linkdiv-dash"> — </span><span class="desc">The triangles show you your currently running apps.</span></a></div>
</div></div></div></div></div>
</div></div>
<div id="launcher-customizing" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Customize the Launcher</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="shell-apps-favorites.html" title="Change which applications show in the Launcher"><span class="title">Change which applications show in the Launcher</span><span class="linkdiv-dash"> — </span><span class="desc">Add, move, or remove frequently-used program icons on the 
    Launcher.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="unity-launcher-change-autohide.html" title="Auto-hide the Launcher"><span class="title">Auto-hide the Launcher</span><span class="linkdiv-dash"> — </span><span class="desc">Show the <span class="gui">Launcher</span> only when you need it.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="unity-launcher-change-size.html" title="Change the size of icons in the Launcher"><span class="title">Change the size of icons in the Launcher</span><span class="linkdiv-dash"> — </span><span class="desc">Make the icons in the Launcher larger or smaller.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
