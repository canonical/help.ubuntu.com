<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Välkommen till Ubuntu</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Välkommen till Ubuntu</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Ubuntu använder <span class="em">Unity</span>, ett nytt sätt att använda din dator. Unity är utformat för att minimera distraktioner, ge dig mer utrymme att arbeta, och hjälper dig få saker utförda.</p>
<p class="p">Den här guiden ska försöka hjälpa dig besvara dina frågor om hur du använder Unity och ditt Ubuntu-skrivbord. Först ska vi titta på några centrala funktioner i Unity, och hur du kan använda dem.</p>
</div>
<div id="unity-overview" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kom igång med Unity</span></h2></div>
<div class="region">
<div class="contents"><div class="media media-image"><div class="inner"><img src="figures/unity-overview.png" class="media media-block" alt="Skrivbordet Unity"></div></div></div>
<div id="launcher-home-button" class="sect"><div class="inner">
<div class="hgroup"><h3 class="title"><span class="title">Programstartaren</span></h3></div>
<div class="region"><div class="contents">
<div class="media media-image floatstart"><div class="inner"><img src="figures/unity-launcher.png" class="media media-block" alt="Programstartaren"></div></div>
<p class="p"><span class="gui">Programstartaren</span> visas automatiskt när du loggar in på ditt skrivbord, och ger dig snabb åtkomst till programmen du oftast använder.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="unity-launcher-intro.html" title="Använda programstartaren">Läs mer om Startaren.</a></span></p></li></ul></div></div></div>
</div></div>
</div></div>
<div id="the-dash" class="sect"><div class="inner">
<div class="hgroup"><h3 class="title"><span class="title">Snabbstartspanelen</span></h3></div>
<div class="region"><div class="contents">
<p class="p"><span class="gui">Ubuntu-knappen</span> sitter vid skärmens övre vänstra hörn, och är alltid det översta objektet i Startaren. Om du klickar på <span class="gui">Ubuntu-knappen</span> kommer Unity visa upp en ytterligare funktion i skrivbordet, <span class="gui">Snabbstartspanelen</span>.</p>
<div class="media media-image"><div class="inner"><img src="figures/unity-dash.png" class="media media-block" alt="Unitys Snabbstartspanel"></div></div>
<p class="p"><span class="em">Snabbstartspanelen</span> är utformad för att göra det lättare att hitta, öppna, och använda program, filer, musik med mera. Om du till exempel skriver ordet "dokument" i <span class="em">Sökfältet</span> kommer Snabbstartspanelen visa dig vilka program som kan hjälpa dig skriva eller redigera dokument. Den kommer också visa dig relevanta mappar och dokument som du har arbetat med nyligen.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="unity-dash-intro.html" title="Hitta program, filer, musik med mera med Snabbstartspanelen">Läs mer om Snabbstartspanelen.</a></span></p></li></ul></div></div></div>
</div></div>
</div></div>
</div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links ">
<a href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord, program &amp; fönster</a><span class="desc"> — <span class="link"><a href="unity-introduction.html" title="Välkommen till Ubuntu">Introduktion</a></span>, <span class="link"><a href="shell-keyboard-shortcuts.html" title="Användbara tangentbordsgenvägar">kortkommandon</a></span>, <span class="link"><a href="shell-windows.html" title="Fönster och arbetsytor">fönster</a></span>…</span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="about-this-guide.html" title="Om denna handbok">Om denna handbok</a><span class="desc"> — Några tips om hur du använder Ubuntu Skrivbordsguide.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
