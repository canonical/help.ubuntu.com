<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Min dator vill inte starta</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="hardware-problems-graphics.html" title="Skärmproblem">Skärmproblem</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="power.html#problems" title="Problem">Strömproblem</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Min dator vill inte starta</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Det finns ett antal skäl till varför din dator inte startar. Detta ämne ger en snabb översikt över några av de möjliga skälen.</p></div>
<div id="nopower" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Datorn är inte ansluten, batteriet är tomt eller kablar lösa</span></h2></div>
<div class="region"><div class="contents"><p class="p">Säkerställ att datorns strömkablar är ordentligt anslutna och att strömkontakterna på slagna. Försäkra dig om att skärmen är ansluten och påslagen också. Om du har en bärbar dator koppla i laddningskabeln (om den har fått slut på batteri). Det kan också vara bra att kontrollera att batteriet är isatt ordentligt (kontrollera undersidan på den bärbara datorn) om det är löstagbart.</p></div></div>
</div></div>
<div id="hardwareproblem" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Problem med datorhårdvaran</span></h2></div>
<div class="region"><div class="contents"><p class="p">En komponent i din dator kan vara trasig eller inte fungera ordentligt. Om detta är fallet kommer du att behöva få din dator reparerad. Vanliga fel omfattar ett trasigt strömaggregat, fel isatta komponenter (som exempelvis minne eller RAM) eller ett trasigt moderkort.</p></div></div>
</div></div>
<div id="beeps" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Datorn piper och stänger sedan av</span></h2></div>
<div class="region"><div class="contents"><p class="p">Om datorn piper flera gånger när du startar den och sedan stänger av sig (eller misslyckas med att starta), kan det vara en indikator på att den har detekterat ett problem. Dessa pip refereras ibland till som <span class="em">pipkoder</span> och mönstret av pip är avsedda att berätta för dig vad felet med datorn är. Olika tillverkare använder olika pipkoder så du måste konsultera manualen för din dators moderkort eller lämna in din dator för reparation.</p></div></div>
</div></div>
<div id="fans" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Datorns fläktar snurrar men ingenting visas på skärmen</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Det första du bör kontrollera är om din skärm är ansluten och påslagen.</p>
<p class="p">Detta problem kan också inträffa på grund av hårdvarufel. Fläktarna kan slås på när du trycker på strömknappen men andra väsentliga delar av datorn kan ha misslyckats att starta. I detta fallet, lämna in din dator för reparation.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="hardware-problems-graphics.html" title="Skärmproblem">Skärmproblem</a><span class="desc"> — Felsök skärm- och grafikproblem.</span>
</li>
<li class="links ">
<a href="power.html#problems" title="Problem">Strömproblem</a><span class="desc"> — Felsök problem med ström och batterier.</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
