<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Öppna program för enheter eller diskar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#removable" title="Flyttbara enheter och externa diskar">Flyttbara enheter och externa diskar</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#photos" title="Foton och digitalkameror">Foton</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#videos" title="Videor och videokameror">Videor</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Öppna program för enheter eller diskar</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan få ett program att starta automatiskt när du ansluter en enhet eller matar in en disk eller ett mediakort. Du vill kanske till exempel att din fotohanterare ska starta när du ansluter en digitalkamera. Du kan också stänga av detta så att ingenting händer när du ansluter något.</p>
<p class="p">För att bestämma vilka program som ska starta när du ansluter olika enheter:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Justeringsverktyg</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Detaljer</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Flyttbar media</span>.</p></li>
<li class="steps">
<p class="p">Hitta din önskade enhet eller mediatyp och välj sedan ett program eller åtgärd för den mediatypen. Se nedan för en beskrivning av de olika typerna av enheter och media.</p>
<p class="p">Istället för att starta ett program kan du också ställa in det så att enheten visas i filhanteraren med alternativet <span class="gui">Öppna mapp</span>. När det händer kommer du att bli tillfrågad vad du vill göra annars kommer inget att hända automatiskt.</p>
</li>
<li class="steps"><p class="p">Om du inte hittar enheten eller mediatypen som du vill ändra i listan (som till exempel Blu-ray-skivor eller eboksläsare) så klicka på <span class="gui">Övriga media…</span> för att se en mer detaljerad lista av enheter. Välj typen av enhet eller media från rullgardinsmenyn <span class="gui">Typ</span> och programmet eller åtgärden i rullgardinsmenyn <span class="gui">Åtgärd</span>.</p></li>
</ol></div></div></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du inte vill att något program ska öppnas automatiskt oavsett vad du ansluter så välj <span class="gui">Fråga aldrig eller starta program när media matas in</span> längst ner i fönstret <span class="gui">Detaljer</span>.</p></div></div></div></div>
</div>
<div id="files-types-of-devices" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Typer av enheter och media</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Ljudskivor</dt>
<dd class="terms"><p class="p">Välj ditt önskade musikprogram eller extraherare för CD-ljud för att hantera ljud-cd. Om du använder dvd (DVD-A) så kan du välja hur de ska öppnas under <span class="gui">Övriga media…</span>. Om du öppnar en ljudskiva med filhanteraren kommer spåren att visas som WAV-filer som du kan spela i vilket musikspelarprogram som helst.</p></dd>
<dt class="terms">Videoskivor</dt>
<dd class="terms"><p class="p">Välj ditt önskade videoprogram för att hantera video-dvd. Använd knappen <span class="gui">Övriga media…</span> för att ställa in ett program för Blu-ray, HD DVD, video-cd (VCD) och super video cd (SVCD). Om dvder eller andra videoskivor inte fungerar korrekt när du matar in dem, se <span class="link"><a href="video-dvd.html" title="Varför spelas inte dvd-filmer upp?">Varför spelas inte dvd-filmer upp?</a></span>.</p></dd>
<dt class="terms">Tomma skivor</dt>
<dd class="terms"><p class="p">Använd knappen <span class="gui">Övriga media…</span> för att välja ett program som skriver skivor för tomma cd, dvder, Blu-ray-skivor och tomma HD-DVD:er.</p></dd>
<dt class="terms">Kameror och foton</dt>
<dd class="terms">
<p class="p">Använd rullgardinsmenyn <span class="gui">Foton</span> för att välja ett fotohanteringsprogram som körs när du ansluter din digitalkamera eller när du matar in ett mediakort från en kamera, exempelvis ett CF-, SD-, MMC- eller MS-kort. Du kan också bara bläddra bland dina foton med hjälp av filhanteraren.</p>
<p class="p">Under <span class="gui">Övriga media…</span> kan du välja ett program för att öppna Kodak-bild-cd, till exempel de som har gjort i en affär. Dessa är vanliga data-cd med JPEG-bilder i en mapp kallad <span class="file">Pictures</span>.</p>
</dd>
<dt class="terms">Musikspelare</dt>
<dd class="terms"><p class="p">Använd ett program för att hantera musikbiblioteket på din bärbara musikspelare eller hantera filerna själv via filhanteraren.</p></dd>
<dt class="terms">E-bokläsare</dt>
<dd class="terms"><p class="p">Använd knappen <span class="gui">Övriga media…</span> för att välja ett program för att hantera böckerna på din e-bokläsare, eller hantera filerna själv via filhanteraren.</p></dd>
<dt class="terms">Programvara</dt>
<dd class="terms">
<p class="p">Vissa skivor och flyttbara media innehåller programvara som är tänkt att köras automatiskt när mediat matas in. Använd alternativet <span class="gui">Programvara</span> för att styra vad som ska hända när media med automatiskt startande program matas in. Du kommer alltid att bli tillfrågad om en bekräftelse innan programvaran körs.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">Kör aldrig program från media du inte litar på.</p></div></div></div></div>
</dd>
</dl></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="files.html#removable" title="Flyttbara enheter och externa diskar">Flyttbara enheter och externa diskar</a></li>
<li class="links "><a href="media.html#photos" title="Foton och digitalkameror">Foton</a></li>
<li class="links "><a href="media.html#music" title="Musik och bärbara ljudspelare">Musik och spelare</a></li>
<li class="links "><a href="media.html#videos" title="Videor och videokameror">Videor</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
