<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Internet verkar vara långsamt</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 19.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk, webb &amp; e-post</a> » <a class="trail" href="net-problem.html.sv" title="Nätverksproblem">Nätverksproblem</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Internet verkar vara långsamt</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Om du använder internet och det verkar långsamt då finns det ett antal saker som kan orsaka att det går långsamt.</p>
<p class="p">Prova att stänga din webbläsare och sedan öppna den igen, samt att prova att koppla ner från internet och sedan ansluta igen. (Att göra detta återställer en massa saker som kan orsaka att internet går långsamt.)</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list">
<p class="p"><span class="em-bold em">En hektisk tid på dagen</span></p>
<p class="p">Internetleverantörer tillhandahåller ställer ofta in internetanslutningar så att de delas mellan flera hushåll. Även om ni ansluter separat via era egna telefonlinjer eller kabelanslutningar, så är anslutningen till resten av internet vid telestationen antagligen delad. Om detta är fallet och många av dina grannar använder internet samtidigt som du kan du uppleva att det går långsamt. Du löper störst risk att uppleva detta vid tidpunkter när dina grannar antagligen använder internet (exempelvis på kvällar).</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Hämta många saker samtidigt</span></p>
<p class="p">Om du eller någon annan som använder din internetanslutning hämtar ner många filer samtidigt eller tittar på videor, så kanske internetanslutningen inte är snabb nog för att hinna med efterfrågan. Om detta är fallet kommer det att upplevas långsammare.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Otillförlitlig anslutning</span></p>
<p class="p">Vissa internetanslutningar är helt enkelt otillförlitliga, speciellt tillfälliga sådana eller de på platser där efterfrågan är stor. Om du är på ett hektiskt café eller på ett konferenscenter så kanske internetanslutningen är allt för upptagen eller helt enkelt otillförlitlig.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Låg signalstyrka för trådlösa anslutningar</span></p>
<p class="p">Om du är trådlöst ansluten till internet (wifi), kontrollera nätverksikonen i systemraden för att se om du har bra trådlös signalmottagning. Om inte kan internet upplevas långsamt för att du inte har en särskilt stark signal.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Att använda en långsammare, mobil internetanslutning</span></p>
<p class="p">Om du har en mobil internetanslutning och märker att den är långsam kan du ha förflyttat dig in i ett område där signalmottagningen är dålig. När detta händer kommer internetanslutningen automatiskt att växla från en snabb ”mobilt bredbands”-anslutning som 3G till en mer tillförlitlig, men långsammare, anslutning som GPRS.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Webbläsaren har problem</span></p>
<p class="p">Ibland inträffar problem som gör webbläsare långsamma. Detta hända på grund av ett antal olika skäl — du kan ha besökt en webbplats som webbläsaren kämpade med att ladda, eller så kan du till exempel ha haft webbläsaren öppen länge. Prova att stänga alla webbläsarens fönster och sedan öppna webbläsaren igen för att se om detta gör någon skillnad.</p>
</li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-problem.html.sv" title="Nätverksproblem">Nätverksproblem</a><span class="desc"> — <span class="link"><a href="net-wireless-troubleshooting.html.sv" title="Felsökning av trådlösa nätverk">Felsök trådlösa anslutningar</a></span>, <span class="link"><a href="net-wireless-find.html.sv" title="Jag kan inte se mitt trådlösa nätverk i listan">hitta ditt trådlösa nätverk</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
