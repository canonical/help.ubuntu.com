<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Hantera program &amp; inställningar via menypanelen</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Hantera program &amp; inställningar via menypanelen</span></h1></div>
<div class="region">
<div class="contents"><p class="p"><span class="gui">Menyfältet</span> är det mörka bandet längst upp i skärmen. Det innehåller fönsterhanteringsknapparna, programmens menyer, och statusmenyerna.</p></div>
<div id="window-management" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Fönsterhanteringsknappar</span></h2></div>
<div class="region">
<div class="contents"><p class="p"><span class="gui">Fönsterhanteringsknapparna</span> visas i fönstrens övre vänstra hörn. I maximerat läge kommer knapparna finnas i skärmens övre vänstra hörn. Klicka på knapparna för att stänga, minimera, maximera, eller återställa fönster.</p></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="shell-windows-states.html" title="Fönsteråtgärder">Fönsteråtgärder</a><span class="desc"> — Återställa, ändra storlek, ordna och dölj.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="app-menus" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Programmenyer</span></h2></div>
<div class="region"><div class="contents">
<p class="p"><span class="gui">Programmenyerna</span> visas som standard till höger om fönsterhanteringsknapparna. Unity döljer programmenyerna och fönsterplaceringsknapparna tills du flyttar din muspekare till skärmens övre vänstra del, eller trycker <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F10</kbd></span></span>. Den här funktionen låter dig se mer av det du jobbar med vid ett givet tillfälle, vilket är särskilt välkommet på mindre skärmar som hos en netbook.</p>
<p class="p">Om du vill kan du ändra det förvalda beteendet, och få dina menyer att sitta tillsammans med fönstrets namnlist för respektive program istället för på menyfältet, samt ange att menyerna alltid skall visas oberoende av musmarkörens position.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="em">Systemmenyn</span> <span class="media"><span class="media media-image"><img src="figures/system-devices-panel.svg" class="media media-inline" alt="Kugghjulsikon"></span></span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">I avsnittet Personligt, klicka på <span class="gui">Utseende</span> och välj fliken <span class="gui">Beteende</span>.</p></li>
<li class="steps"><p class="p">Under <span class="gui">Visa menyerna för ett fönster</span>, välj <span class="gui">I fönstrets namnlist</span>.</p></li>
<li class="steps"><p class="p">Under <span class="gui">Menyernas synlighet</span>, välj <span class="gui">Visas alltid</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="status-menus" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Statusmenyer</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Ubuntu har flera olika <span class="gui">statusmenyer</span> (ibland kallade <span class="gui">indikatorer</span>) till höger på menyfältet. Statusmenyerna är en bekvämt belägen plats där du kan kontrollera och ändra tillståndet för din dator och dina program.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Vissa av ikonerna som används av indikatormenyerna ändras med programmets status.</p></div></div></div></div>
<p class="p">Andra program, som <span class="app">Tomboy</span> eller <span class="app">Transmission</span>, kan också lägga till indikatormenyer på panelen.</p>
<div class="list ui-expander">
<div class="yelp-data yelp-data-ui-expander" dir="ltr" data-yelp-expanded="false"></div>
<div class="inner">
<div class="title title-list"><h3><span class="title">Lista över statusmenyer och vad de gör</span></h3></div>
<div class="region"><ul class="list" style="list-style-type:disc">
<li class="list">
<p class="p"><span class="em">Nätverksmeny</span> <span class="media"><span class="media media-image"><img src="figures/network-offline.svg" class="media media-inline" alt="Frånkopplad nätverksikon"></span></span></p>
<p class="p">Anslut till <span class="link"><a href="net-wired-connect.html" title="Anslut till ett trådbundet (Ethernet) nätverk">trådbundna</a></span>, <span class="link"><a href="net-wireless-connect.html" title="Anslut till ett trådlöst nätverk">trådlösa</a></span>, <span class="link"><a href="net-mobile.html" title="Anslut till mobilt bredband">mobila</a></span>, och <span class="link"><a href="net-vpn-connect.html" title="Anslut till ett VPN">VPN-</a></span>nätverk.</p>
</li>
<li class="list">
<p class="p"><span class="em">Meny för inmatningskällor</span> <span class="media"><span class="media media-image"><img src="figures/indicator-keyboard-En.svg" class="media media-inline" alt="Ikon för inmatningskällor"></span></span></p>
<p class="p">Välj tangentbordslayout/indatakälla, <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">anpassa indatakällor</a></span>.</p>
</li>
<li class="list">
<p class="p"><span class="em">Bluetooth-meny</span> <span class="media"><span class="media media-image"><img src="figures/bluetooth-active.svg" class="media media-inline" alt="Bluetooth-ikon"></span></span></p>
<p class="p">Skicka eller ta emot filer via <span class="link"><a href="bluetooth.html" title="Bluetooth">Bluetooth</a></span>. Den här menyn är dold när ingen Bluetooth-enhet upptäcks och stöds.</p>
</li>
<li class="list">
<p class="p"><span class="em">Meddelandemeny</span> <span class="media"><span class="media media-image"><img src="figures/indicator-messages.svg" class="media media-inline" alt="Meddelandeikon"></span></span></p>
<p class="p">Starta och ta enkelt emot inkommande aviseringar från meddelandeprogram, inklusive e-post, sociala nätverk, och internet-chat.</p>
</li>
<li class="list">
<p class="p"><span class="em">Batterimeny</span> <span class="media"><span class="media media-image"><img src="figures/battery-100.svg" class="media media-inline" alt="Batteri-ikon"></span></span></p>
<p class="p">Kontrollera din bärbara dators laddning. Den här menyn är dold när inget batteri upptäcks.</p>
</li>
<li class="list">
<p class="p"><span class="em">Ljudmeny</span> <span class="media"><span class="media media-image"><img src="figures/audio-volume-high-panel.svg" class="media media-inline" alt="Ljudikon"></span></span></p>
<p class="p">Ställ in <span class="link"><a href="sound-volume.html" title="Ändra ljudvolymen">volym</a></span>, anpassa <span class="link"><a href="media.html" title="Ljud, video och bilder">ljudinställningar</a></span>, och styr mediaspelare som <span class="app">Rhythmbox</span>.</p>
</li>
<li class="list">
<p class="p"><span class="em">Klocka</span></p>
<p class="p">Kom åt aktuell tid och datum. Möten från <span class="link"><a href="clock-calendar.html" title="Kalendermöten">Kalender</a></span>-programmet kan också visas här.</p>
</li>
<li class="list">
<p class="p"><span class="em">Systemmeny</span> <span class="media"><span class="media media-image"><img src="figures/system-devices-panel.svg" class="media media-inline" alt="Kugghjulsikon"></span></span></p>
<p class="p">Kom åt detaljinformation om din dator, den här hjälpen, och <span class="link"><a href="prefs.html" title="Inställningar för användare och system">systeminställningar</a></span>. Växla användare, lås skärmen, logga ut, gå i vänteläge, starta om, eller stäng av din dator.</p>
</li>
</ul></div>
</div>
</div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="index.html" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li>
<li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
