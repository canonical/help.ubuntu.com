�PNG

   IHDR  v      tYf   �zTXtRaw profile type exif  x�mPm� ��)vT8�]�d7���I��%>��'�����#'.M�֊V��������V�"z�C�є-�%��N�V<�����$$�Hlׄr�ˏP<D>Q6g!!�3�B�ǤU����x��N[������Ͷ�{�r>HI����P7����V�6.�&�E��i��"Z�/a  �iCCPICC profile  x�}�=H�@�_S�"�q�P����U(B�P+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�F�iV�,�鶙N&�lnU�"�D0Qf�1'I)���{�z�Y���}j�b@@$�e�ioOo��}�(+�*�9�I$~�����ό���<q�X,v����dj�S�1U�)_�z�r��Uj�uO��p^_Y�:�a$��%H���2*��U'�B��>�!�/�K!W��B������w�Var�K
'����B�@��8�ǎ�<������W��'���;����붦��;���!��+i
��~Fߔ"�@��[k�@��J� ��h���}����ۿgZ�� ��r�(˞�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:47ac6055-f470-439b-91da-30d907781218"
   xmpMM:InstanceID="xmp.iid:c0d485b8-178f-4d2b-a158-862b6640abd2"
   xmpMM:OriginalDocumentID="xmp.did:be77ea3a-9017-43bb-aad0-4a19e1ee86cc"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679601894936326"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T21:04:54+01:00"
   xmp:ModifyDate="2023:03:23T21:04:54+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:1254538a-f7c7-48b1-a42a-867169133b6e"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T21:04:54+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>:�C   	pHYs  �  ��+   tIME�	:��   tEXtComment Created with GIMPW�  MIDATx��yp[�}���~8 o��%�,'�!��S;n��$v��NƝ$Mf��t�?�_;�N�i&m���I\'>#Y�m)�-�K�n��D�& �$�w����H��R	����<<������������`0��e&�,��`07(��W$�&�X<fۄ�/�B�,�BA���&$�H�R�f!�N�M<���4�! �l6��r9� �ec
#���B!��X~0e��g�vJ!�g��,����Ü��$��1�ѓ�TUU5��,W��&�ɱ��ښ ���i���a�Y�0�`�f8EQQ L�'�9���%�����Yn�?�d2���ƭN��8���������9�9������999��9����M�W���  �e��$���1���i������1�	� �`[V�Zt]�8��8f0�9B,��uXHٓH&?س7�H��y���kn��7���j �P�L#D(-�$��&i��.i@�N' ��`*���|��F��p8�7�B�I)]��`Ș4oQæQ�C��$c&L,�(s�����̯FP*I��4PT���Z��8�癊ɘIPJ)�/oN�<����u�4M�ӤE�&{J�������45a�Bz6;2:j�<��$��*���Y��dzdd��[>�PU�ꪐ�( BE'&"��. !��Y]*v��L�����F�k� H�i:OMJ�&���:q,:6��|}c���w{������E��w~�0m*�Y�E�@.�*'�i�;op�i>K5��u;Z����r��iǂ��j�ɰj�H�mԌw���;�H
V����'�N;��=縢(~���E���K��7� et��% ������
1�ҩt	�K �f�ɏZp��T�E�R:99i�6����M���7��z��Xt"��?��Z��5BM�7,z����k����u�c�[k*�}2+���>�rg�|��^��W�OJ(� _8o=�"��n�Q�)��{`���^i�v
 X�S����96��Ώ4Y�O���b)%�J����"�,٬��~�)-���%}5|Q��b�|��޾K3�޼q���s��Rt������E_�ſ���ɏ��F*�6 $'�C'�_��rtl��1Y-�<b�)S�g+Y�0A-B+�>k"k=������ ����ɬ��j�$����yMaƝ7\K�Nd��n���xL	6�x�A��y6K�F��&ђ��R��ܘ�I)��k�_��9�F愘�`S�H�v��^7��g�9��=<�6v8������{� S1�'��B)<���E��i,����X*�5D�)�T��gb$,�s��]��<T;��:2�Έ�r�<�Ek����ۥI�<J.��ӯkbZVǪ��=��s�>[[[c��Bś��*B�t9�'{��Es�őݹ/��+��s�CA���'?~+<�)��CCw�|���{�����"���C���ԡ�]z6��S�+�M.mR�� )�ưi.g �r+�G�V�0)"xV�:w���� �R��1�mX',�X4����5^���U{��7|�����j�x�*��P<�д�Sg���yBȹ��GF�\��ԩ\.w���˗Ñ{Re�Xث�_K"�ѥRP�.�[����ƅ^��i��]���o>��7�o��_�V
��w<��_�>��v�:�����/w��?D�o��+4os�	kW�A�t���"�������R2�*|<����o���3���B���N]י�-g��O���]��}.�C�NQj��|]W�9���3W����o�mٶ(
׺�G�;{z��#��b�K1y#���L��f��m�zƲ���IJIa��ɖi�����r���~z��C��:��'�7b�������U�%e�r-a�S���--Kxה�H��q�d*��z�~�s ��۷c�. ��/�29#1~y��*p" �����l�r�m�;w�t�ϗz��q�����y�����ڝ��7_�JF��^��p�@�ȱ�7n�z�t{k�����A��ް~�W�H����htttl����IY�R�k����_?���ߞ�� 0)����5��W��������i����$�ɺ�ڕ��]����沊�t=��4A�������y��5�$�8�-I�Dl⾭[��e�K-�"O-�&�2B BaV ��x�l~�OFFG��8��G�4���x���q{[�V4�"�J���qwW[� gϝ'�Z���ڪ�ݖm���&��p$R
@,�tY����Jȥ�~�4}^_}]-{�%�N���A�0�\R牖膧�zj9�����O��'?��W�:�c|����?��O���+W�����"W_�P��1QDX@X��9�����xeehd�*W��g��ukք#�����A����z)зw�,��ٻohx�ͷ��p88�C����]/To���MlV�ʲ�Sz��辻��'WN 2s�ݱZ���{��t��+��?�} B�� 
;���w�r4}��W�ɔ�(�,��nEQ����߻W�C��t= ���}��'��]e$bN9��-���`"�0�~Ma��v����yx��`   �T ���w(>m�G���8t�H6�۳�C˲��m���3{z$I�'������C۶��N��N�R;w�N�R<���R�a�;K8�g�j���h�h��"����m���׭������@}�Ux��	�"�*��[�s���n�ro>�?���מ�N�,:<n�5��kA6mX���H4��C��_��4!$�H�Z�rfK!J��7�\�ѱ~�Z&aަ`@.^�G (B�iJ9ĭ���?�vs.�I��h"�TE�5�;ɤ��i��[u�]�>�� 'Nt��4����mjl�v��5�5;v��v�}<�?��_�}>���8\�q٬�FJ�7wС�ÿˉ���=�r�R�8�=�*
Bh`p(rWW[�����'gΙ��z���ZZ0Ɨ�����]���*<x�K���z{��@��2� @$���z�J�0����jk��sk��V�d0�i\��,Q=~M  ���'_���_������u�=a�*U5�<�, ڦ��=������6��� c���xǆ�~�������.Z�]_W7spf�)����מ�8�ͷ��9AӴ�Q�f*f�ʘ��S+{_����0���?_���7eBڂ�lo[ӱ�;M�G"��{/��o&4˶_�<�qLj*{ij���YVdY�$Y��'��<�������8��r]eʲ���_8s��Ş�4=:J����B�Pd���l��[�ĒPj���n�|Ss�7o����%t,��V1�P�[~R�M��-�b����P��SݧN�~����.\�C�wJ�-n�wۇG��l�����������}0X$ ��N\�ZZ[�����������Ӆ8 !Դ�q�w��IF�'3��������Ԡ+���/>�1�����e1�{�������<�&���j��K/ȭ��mm�P�#�ꬪ5�m.0����/<�H�����-�D"QA�y��VVV�:}fl|����̹s]G�~�ٹe�&�Xn;sA?�OP � �h@<�1�`�m˶m�^hwZ�����=p����`8�-�V���r�\�uu�T��t(��qW��%���n����/^��
(�u��t8T���]�����j����
�&�EU��)���oϜ=��{��`�d&�z��͛6.���d�/t	���P��9�QN���W?lo�V�$��Qaΰ���^M=���55�����x�����**��� �$��55�-�щ	۶ׯ]���ÑHǪ��Vɲ\WS�p8V46�lo�'�ա����ˇD<��h 09��e��'1(��ß����df�Bb|(>ty{���7?�i}������"��_9�9�h��4%h	B0�4mEcc6�min�eyb"���������]�`0�
��DB���f��;<<�Ըbúu�I�TW[ì�|�d2"?�X���󅍆ߺTq��b� ��!ba,�mJ)!��D�xJI����^���� ����hlBUԆ��P0XYYO$�~_ӊ�d25��h���r*�Tr�PU��_����H$�V����r:�u��DB׳��r:UU���:��k!!���r����饔�9�%IR�-���7����H$�q�z�����lI;�á��e���T�0��$��ݢ ض��x>�ۥ�����!2��EÅw#�c>�,���82zՊq΅�-���p� �L�l��m�O����+�v}|��{O>��~���)���7wD��O|�5�ͫ�jZ|���ù|�Ҋ�z koqk$�s<� QuIn?vV^>{̚����D,ӶI�t<�+N��w0Ŏ�ԙ3���<?���_[���# :-"B�i� �z�d�&l�;B�eY����Yn�9［��z��9��n��أ�����ٳ/~���$+�h4�(͝*+�~_>�E�$EN�ӥI���ơ��������w)_�趥�	cdM��H��UU7�d(�[F�s�vmm�W_h]����ݻ;8S����X��o��U��@�&�ޥe";,|�W݀9J5�"8<��6��~
��݈yA�\~̳���Rf2ͳ������S��|���8��\.o*�c��7�U~���E�V~(I�ϸ��%�BM���( `\¤* *tޠR�ۙ�ޢ���D��y��]s�|����׺��B[喍�֌�'��,���t6T�+��!�8֩�LꂅM�j��!��'* ��<��ۜc�Xgz�wz{���ϫg�� in��cY֎�Q>�|ޞ޾H$�iWM܌�b�T�'gY���
�q9���^�kI��%6
(!M��rs�	�
�*I%�E�RB}^Ot"FnqOB��trGlk�$�3���Ng,��r7�ۖElK�g/5V��A� T*uM�j��0߿�*���� �Թ�1Ye���#LZg��+�($
HdJ6s)t�ca�-�W����/^���{��8���ݽi#F(5C������RJ�i�6i�"+�MM�)ĶIj[������4Iۖe[�LI�gJ���~�Ӽ�v�(������K�<�N�L�{�i@�S�s	˪2���,�$��dR�$6��1�0���ˡ�EQ�|�DE�}��۲T���&��p<p�}�t�4�[=��Ü��t9��dlb�|�4��:3�ǲ-B*]�dF��,�&vi�&�PPOg�����MO&���D��0��!Pd���bJJi2�N�&)���9������`�a�b�|>ǌ�1ױ`�*l�>�Q~e3rBL��`0ƲV
>�����`0�M�� �r��Yt�    IEND�B`�