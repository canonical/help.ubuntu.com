<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Control Groups</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="lxc.html" title="LXC">Föregående</a><a class="nextlinks-next" href="cgroups-overview.html" title="Översikt">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Control Groups</h1></div>
<div class="region">
<div class="contents">
<p class="para">
Control groups (cgroups) are a kernel mechanism for grouping, tracking,
and limiting the resource usage of tasks.  The kernel-provided administration
interface is through a virtual filesystem.  Higher level cgroup
administration tools have been developed, including libcgroup and
lmctfy.  Additionally, there is guidance at freedesktop.org
for how applications can best cooperate using the cgroup filesystem
interface (see Resources).
  </p>
<p class="para">
As of Ubuntu 14.04, the cgroup manager (cgmanager) is available as
another cgroup administion interface.  It's goal is to respond to dbus
requests from any user, allowing him to administer only those cgroups
which have been delegated to him.
  </p>
<p class="para">
<a class="xref" href="cgroups-overview.html" title="Översikt">Översikt</a> will describe cgroups in more detail.
<a class="xref" href="cgroups-fs.html" title="Filesystem">Filesystem</a> will describe the long-standing cgroups filesystem
interface.  <a class="xref" href="cgroups-manager.html" title="Manager">Manager</a> will describe the cgroup
manager.
  </p>
</div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="cgroups-overview.html" title="Översikt">Översikt</a></li>
<li class="links"><a class="xref" href="cgroups-fs.html" title="Filesystem">Filesystem</a></li>
<li class="links"><a class="xref" href="cgroups-delegation.html" title="Delegation">Delegation</a></li>
<li class="links"><a class="xref" href="cgroups-manager.html" title="Manager">Manager</a></li>
<li class="links"><a class="xref" href="cgroups-resources.html" title="Resurser">Resurser</a></li>
</ul></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="lxc.html" title="LXC">Föregående</a><a class="nextlinks-next" href="cgroups-overview.html" title="Översikt">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
