<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Filegenskaper</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Filegenskaper</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">För att visa information om en fil eller mapp, högerklicka på den och välj <span class="gui">Egenskaper</span>. Du kan också markera filen och trycka <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Retur</kbd></span></span>.</p>
<p class="p">Filegenskapsfönstret visar information om filtyp, filstorlek, och när du senast ändrade den. Om du behöver den här information ofta kan du visa den i <span class="link"><a href="nautilus-list.html" title="Inställningar för filhanterarens listkolumner">listvyns kolumner</a></span> eller <span class="link"><a href="nautilus-display.html#icon-captions" title="Ikontext">ikontext</a></span>.</p>
<p class="p">Information som visas i fliken <span class="gui">Grundläggande</span> förklaras nedanför. Det finns också flikar för <span class="gui"><span class="link"><a href="nautilus-file-properties-permissions.html" title="Ange filrättigheter">Rättigheter</a></span></span> och <span class="gui"><span class="link"><a href="files-open.html#default" title="Ändra förvalt program">Öppna med</a></span></span>. För vissa filtyper, som bilder och videor, finns en ytterligare flik som visar information om dimensioner, längd, och kodek.</p>
</div>
<div id="basic" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Grundläggande egenskaper</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms"><span class="gui">Namn</span></dt>
<dd class="terms"><p class="p">Du kan döpa om filen genom att ändra i det här fältet. Du kan också döpa om en fil utanför egenskapsfönstret. Se <span class="link"><a href="files-rename.html" title="Byt namn på en fil eller mapp">Byt namn på en fil eller mapp</a></span>.</p></dd>
<dt class="terms"><span class="gui">Typ</span></dt>
<dd class="terms">
<p class="p">Detta hjälper dig identifiera filens typ, som PDF-dokument, OpenDocument-text, eller JPEG-bild. Filtypen avgör bland annat vilka program som kan öppna filen. Se <span class="link"><a href="files-open.html" title="Öppna filer med andra program">Öppna filer med andra program</a></span> för ytterligare information.</p>
<p class="p">Filens <span class="em">MIME-typ</span> visas i parenteser; MIME-typ är en standardmetod som datorer använder för att hänvisa till filtypen.</p>
</dd>
<dt class="terms">Innehåll</dt>
<dd class="terms"><p class="p">Det här fältet visas om du tittar på egenskaperna för en mapp istället för en fil. Det hjälper dig att se antal objekt i mappen. Om mappen innehåller andra mappar kommer varje underliggande mapp räknas som ett objekt, även om det innehåller andra objekt. Varje fil räknas också som ett objekt. Om mappen är tom kommer Innehåll visa <span class="gui">tom</span>.</p></dd>
<dt class="terms">Storlek</dt>
<dd class="terms">
<p class="p">Det här fältet visas om du tittar på en fil (inte en mapp). Filstorleken visar dig hur mycket diskutrymme den tar upp. Detta är också en indikator för hur länge det kommer ta att ladda ner en fil eller skicka den med e-post (stora filer tar lång tid att skicka/ta emot).</p>
<p class="p">Storlekar kan anges i byte, KB, MK, eller GB; för de tre sista kommer storlek i byte också visas i parenteser. Tekniskt sett är 1 KB 1024 byte, 1 MB är 1024 KB, och så vidare.</p>
</dd>
<dt class="terms">Plats</dt>
<dd class="terms"><p class="p">Platsen för varje fil på din dator anges som dess <span class="em">absoluta sökväg</span>. Detta är en unik "adress" för filen på din dator, bestående av en lista av de mappar du skulle behöva navigera genom för att hitta filen. Om till exempel Jim har en fil som heter <span class="file">Resume.pdf</span> i sin Hemmapp skulle dess plats vara <span class="file">/home/jim/Resume.pdf</span>.</p></dd>
<dt class="terms">Volym</dt>
<dd class="terms"><p class="p">Filsystemet eller enheten som filen lagras på. Detta visar dig var filen fysiskt lagras, till exempel på en hårddisk eller en CD, eller en <span class="link"><a href="nautilus-connect.html" title="Bläddra bland filer på en server eller nätverksdelning">nätverksdelning eller filserver</a></span>. Hårddiskar kan delas upp i flera <span class="link"><a href="disk-partitions.html" title="Hantera volymer och partitioner">diskpartitioner</a></span>; partitionsnamnet kommer också visas under <span class="gui">Volym</span>.</p></dd>
<dt class="terms">Ledigt utrymme</dt>
<dd class="terms"><p class="p">Detta visas bara för mappar. Det visar hur mycket diskutrymme som finns tillgängligt på disken som mappen finns på. Detta gör det lättare att se om hårddisken är full.</p></dd>
<dt class="terms">Åtkommen</dt>
<dd class="terms"><p class="p">Tid och datum då filen senast öppnades.</p></dd>
<dt class="terms">Ändrad</dt>
<dd class="terms"><p class="p">Tid och datum när filen senast ändrades och sparades.</p></dd>
</dl></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="nautilus-file-properties-permissions.html" title="Ange filrättigheter">Ange filrättigheter</a><span class="desc"> — Styr vem som kan visa och redigera dina filer och mappar.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
