<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Min dator blir väldigt varm</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="power.html#problems" title="Problem">Strömproblem</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Min dator blir väldigt varm</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">De flesta datorer blir varma efter ett tag och visa kan blir riktigt varma. Detta är normalt: det är helt enkelt en del av sättet på vilket datorn kyler sig själv. Om datorn blir allt för varm kan det vara ett tecken på att den överhettas, vilket potentiellt kan orsaka skador.</p>
<p class="p">De flesta bärbara datorer blir ganska varma när du använt dem ett tag. Det är vanligtvis inget att oroa sig för — datorer producerar mycket värme och bärbara datorer är väldigt kompakta så de måste avge sin värme snabbt och deras ytterhölje värms upp som ett resultat. Vissa bärbara datorer blir dock för varma och kan bli obehagliga att använda. Detta är normalt ett resultat av dåligt designade kylsystem. Du kan ibland köpa extra kylningstillbehör som täcker botten på den bärbara datorn och ger en mer effektiv kylning.</p>
<p class="p">Om du har en stationär dator som känns varm vid beröring kan den ha otillräcklig kylning. Om detta bekymrar dig kan du köpa extra kylningsfläktar eller kontrollera att kylningsfläktarna och ventilationen inte är blockerade av damm eller något annat. Det kan också vara bra att överväga att placera datorn på en bättre ventilerad plats — om den placeras i trånga utrymmen (till exempel i ett skåp) kan det vara så att kylsystemet i datorn inte kan avge värme och cirkulera kall luft snabbt nog.</p>
<p class="p">Vissa personer är bekymrade om hälsoeffekterna av att använda bärbara datorer. Det finns indikationer på att förlängd användning av en varm, bärbar dator i ditt knä möjligt skulle kunna reducera (manlig) fruktbarhet och det finns rapporter om mindre brännmärken (i extrema fall). Om du är bekymrad om dessa potentiella problem kan det vara bra att ta kontakt med en praktiserande läkare för råd. Naturligtvis kan du helt enkelt välja att inte ha den bärbara datorn i ditt knä.</p>
<p class="p">De flesta moderna datorer kommer att stänga ner sig själva om de blir allt för varma, för att förhindra att de själva blir skadad. Om din dator stänger ner sig ofta kan detta vara orsaken. Om din dator överhettas kommer du förmodligen att behöva få den reparerad.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="power.html#problems" title="Problem">Strömproblem</a><span class="desc"> — Felsök problem med ström och batterier.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
