<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Översikt</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="cgroups.html" title="Control Groups">Control Groups</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups.html" title="Control Groups">Föregående</a><a class="nextlinks-next" href="cgroups-fs.html" title="Filesystem">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Översikt</h1></div>
<div class="region"><div class="contents">
<p class="para">
Cgroups are the generalized feature for grouping tasks.  The actual
resource tracking and limits are implemented by subsystems.  A
hierarchy is a set of subsystems mounted together.  For instance,
if the memory and devices subsystems are mounted together under
/sys/fs/cgroups/set1, then any task which is in "/child1" will
be subject to the corresponding limits of both subsystems.
  </p>
<p class="para">
Each set of mounted subsystems consittutes a 'hierarchy'.  With
exceptions, cgroups which are children of "/child1" will be
subject to all limits placed on "/child1", and their resource
usage will be accounted to "/child1".
  </p>
<p class="para">
The existing subsystems include:
  </p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist"><p class="para"><span class="em emphasis">cpusets</span>: fascilitate assigning a set of
CPUS and memory nodes to cgroups.
  Tasks in a cpuset cgroup may only be scheduled on CPUS assigned to that
  cpuset.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> blkio </span>: limits per-cgroup block io.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> cpuacct </span>: provides per-cgroup cpu usage accounting.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> devices </span>: controls the ability of tasks to create or use devices nodes
  using either a blacklist or whitelist.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> freezer </span>: provides a way to 'freeze' and 'thaw' whole cgroups.  Tasks
  in the cgroup will not be scheduled while they are frozen.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> hugetlb </span>: fascilitates limiting hugetlb usage per cgroup.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> memory </span>: allows memory, kernel memory, and swap usage to be tracked
  and limited.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> net_cls </span>: provides an interface for tagging packets based on the
  sender cgroup.  These tags can then be used by tc (traffic controller)
  to assign priorities.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> net_prio </span>: allows setting network traffic priority on a per-cgroup
  basis.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> cpu </span>: enables setting of scheduling preferences on per-cgroup basis.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis"> perf_event </span>: enables per-cpu mode to monitor only threads in certain
  cgroups.</p></li>
</ul></div>
<p class="para">
In addition, named cgroups can be created with no bound
subsystems for the sake of process tracking.  As an example,
systemd does this to track services and user sessions.
  </p>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups.html" title="Control Groups">Föregående</a><a class="nextlinks-next" href="cgroups-fs.html" title="Filesystem">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
