<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Lägg till fler programförråd</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="addremove.html" title="Lägg till &amp; ta bort mjukvara">Lägg till/ta bort program</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Lägg till fler programförråd</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Program kan hämtas från tredjepartskällor, såväl som från Ubuntus standardprogramarkiv. Om du vill installera program från ett tredjepartsarkiv måste du lägga till det till Ubuntus lista över tillgängliga arkiv.</p>
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents">
<p class="p">Lägg bara till programarkiv från källor du litar på!</p>
<p class="p">Externa arkiv kontrolleras inte för säkerhet eller stabilitet av Ubuntumedlemmar, och kan innehålla program som är skadliga för din dator.</p>
</div></div></div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Installera andra arkiv</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ikonen <span class="app">Programcentral för Ubuntu</span> i programstartaren, eller sök efter Programcentral i sökraden i <span class="app">Dash</span>.</p></li>
<li class="steps"><p class="p">När programcentralen startas, klicka på <span class="guiseq"><span class="gui">Redigera</span> ▸ <span class="gui">Programkällor</span></span></p></li>
<li class="steps"><p class="p">Du kommer få skriva in ditt lösenord. När du har gjort det, byt till fliken <span class="gui">Övriga program</span>.</p></li>
<li class="steps">
<p class="p">Klicka på <span class="gui">Lägg till</span> och skriv in APT-raden för arkivet. Detta bör finnas tillgängligt från arkivets webbplats, och bör se ut så här:</p>
<p class="p">
        <span class="code">deb http://archive.ubuntu.com/ubuntu/ trusty main</span>
      </p>
</li>
<li class="steps"><p class="p">Klicka på <span class="gui">Lägg till källa</span> och stäng sedan fönstret Program &amp; uppdateringar. Programcentralen kommer att söka igenom dina programkällor för nya uppdateringar.</p></li>
</ol></div>
</div></div>
</div>
<div id="canonical-partner" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Aktivera förrådet Canonical-partners</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Canonicals partnerarkiv tillhandahåller en del slutna program; de kostar inget, men använder inte öppen källkod. Där finns program som <span class="app">Skype</span>, <span class="app">Adobe Reader</span> och <span class="app">Adobe Flash Plugin</span>. Programmen i det här arkivet kommer visas bland Ubuntus programcentrals sökträffar, men går inte att installera om inte arkivet har aktiverats.</p>
<p class="p">För att aktivera arkivet, följ stegen ovan för att öppna fliken <span class="gui">Övriga program</span> i <span class="app">Program &amp; uppdateringar</span>. Om du ser arkivet <span class="gui">Canonical-partners</span> i listan, se till att det har kryssats för och stäng sedan fönstret Program &amp; uppdateringar. Om du inte ser det, klicka på <span class="gui">Lägg till</span> och skriv in:</p>
<p class="p">
      <span class="code">deb http://archive.canonical.com/ubuntu trusty partner</span>
    </p>
<p class="p">Klicka på <span class="gui">Lägg till källa</span> och stäng sedan fönstret Program &amp; uppdateringar. Vänta en liten stund medan Ubuntus programcentral laddar ner arkivinformationen.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="addremove.html" title="Lägg till &amp; ta bort mjukvara">Lägg till &amp; ta bort mjukvara</a><span class="desc"> — <span class="link"><a href="addremove-install.html" title="Installera fler program">Installera</a></span>, <span class="link"><a href="addremove-remove.html" title="Ta bort ett program">ta bort</a></span>, <span class="link"><a href="addremove-sources.html" title="Lägg till fler programförråd">extra förråd</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="addremove-ppa.html" title="Lägg till ett Privat PaketArkiv (PPA)">Lägg till ett Privat PaketArkiv (PPA)</a><span class="desc"> — Lägg till PPA:er för att hjälpa till att testa experimentell kod eller specialprogram.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
