<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Tangentbordsnavigation</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 19.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="keyboard.html.sv" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 19.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="keyboard.html.sv" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 19.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="a11y.html.sv" title="Hjälpmedel">Hjälpmedel</a> › <a class="trail" href="a11y.html.sv#mobility" title="Rörelsehinder">Rörelsehinder</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Tangentbordsnavigation</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Denna sida beskriver tangentbordsnavigering för personer som inte kan använda en mus eller annat pekdon eller som vill använda tangentbordet så mycket som möjligt. För snabbtangenter som är användbara för alla användare, se <span class="link"><a href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar">Användbara tangentbordsgenvägar</a></span> istället.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du inte kan använda ett pekdon som exempelvis en mus kan du kontrollera musmarkören med hjälp av den numeriska delen på ditt tangentbord. Se <span class="link"><a href="mouse-mousekeys.html.sv" title="Klicka och flytta muspekaren med det numeriska tangentbordet">Klicka och flytta muspekaren med det numeriska tangentbordet</a></span> för detaljer.</p></div></div></div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h2><span class="title">Navigera i användargränssnitt</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td>
<p class="p"><span class="key"><kbd>Tabb</kbd></span> och</p>
<p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p>
</td>
<td>
<p class="p">Flytta tangentbordsfokus mellan olika kontroller. <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span> flyttar mellan grupper av kontroller, som exempelvis från en sidopanel till huvudinnehållet. <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span> kan också bryta loss från en kontroll som själv använder <span class="key"><kbd>Tabb</kbd></span>, till exempel ett textområde.</p>
<p class="p">Håll ner <span class="key"><kbd>Skift</kbd></span> för att flytta fokus i omvänd ordning.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p">Piltangenter</p></td>
<td style="border-top-style: solid;"><p class="p">Flytta markering mellan objekt inom en kontroll, eller mellan en mängd av relaterade kontroller. Använd piltangenterna för att fokusera på knappar i en verktygsfält, markera objekt i en lista eller ikonvy eller markera radioknappar från en grupp.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+Piltangenter</span></p></td>
<td style="border-top-style: solid;"><p class="p">I en list- eller ikonvy, flytta tangentbordsfokus till ett annat objekt utan att ändra vilket objekt som är markerat.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Shift</kbd></span>+Piltangenter</span></p></td>
<td style="border-top-style: solid;">
<p class="p">I en list- eller ikonvy, markera alla objekt från och med det för närvarande valda objektet till och med det nyligen fokuserade objektet.</p>
<p class="p">I en trädvy kan objekt med underordnade objekt expanderas och fällas ihop så att de underordnade objekten visas eller döljs. Expandera genom att trycka <span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>→</kbd></span></span>, fäll ihop genom att trycka <span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>←</kbd></span></span>.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Blanksteg</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Aktivera ett fokuserat objekt som exempelvis en knapp, kryssruta eller listobjekt.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">I en list- eller ikonvy, markera eller avmarkera det fokuserade objektet utan att avmarkera andra objekt.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Alt</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Håll ner <span class="key"><kbd>Alt</kbd></span>-tangenten för att visa <span class="em">snabbtangenter</span>: understrukna bokstäver i menyobjekt, knappar och andra kontroller. Tryck på <span class="key"><kbd>Alt</kbd></span> samt den understrukna bokstaven för att aktivera en kontroll, precis som om du hade klickat på den.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Esc</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Stäng en meny, snabbvalsmeny, växlare eller dialogruta.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>F10</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Öppna den första menyn på menyraden i ett fönster. Använd piltangenterna för att navigera i menyerna.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span>+<span class="key"><kbd>F10</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Öppna programmenyn på systemraden.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;">
<p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>F10</kbd></span></span> eller</p>
<p class="p"><span class="key"><a href="keyboard-key-menu.html.sv" title="Vad är Windows-tangenten?"><kbd>Menu</kbd></a></span></p>
</td>
<td style="border-top-style: solid;"><p class="p">Poppa upp snabbvalsmenyn för den aktuella markeringen som om du hade högerklickat.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>F10</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">I filhanteraren, poppa upp snabbvalsmenyn för den aktuella mappen som om du hade högerklicka på bakgrunden och inte på något objekt.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;">
<p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>PageUp</kbd></span></span></p>
<p class="p">och</p>
<p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>PageDown</kbd></span></span></p>
</td>
<td style="border-top-style: solid;"><p class="p">I ett gränssnitt med flikar, växla till fliken till vänster eller höger.</p></td>
</tr>
</table></div>
</div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h2><span class="title">Navigera skrivbordet</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td>
<p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F1</kbd></span></span> eller</p>
<p class="p">tangenten <span class="key"><a href="keyboard-key-super.html.sv" title="Vad är Super-knappen?"><kbd>Super</kbd></a></span></p>
</td>
<td><p class="p">Växla mellan översiktsvyn <span class="gui">Aktiviteter</span> och skrivbordet. I översiktsvyn kan du börja skriva för att omedelbart söka bland dina program, kontakter och dokument.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-windows-switching.html.sv" title="Växla mellan fönster">Växla snabbt mellan fönster</a></span>. Håll ner <span class="key"><kbd>Skift</kbd></span> för omvänd ordning.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>`</kbd></span></span></p></td>
<td style="border-top-style: solid;">
<p class="p">Växla mellan fönster från samma program, eller från det markerade programmet efter <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span>.</p>
<p class="p">Detta kortkommando använder <span class="key"><kbd>`</kbd></span> på amerikanska tangentbord, där tangenten <span class="key"><kbd>`</kbd></span> sitter ovanför <span class="key"><kbd>Tabb</kbd></span>. På alla andra tangentbord är kortkommandot <span class="key"><kbd>Super</kbd></span> samt tangenten ovanför <span class="key"><kbd>Tabb</kbd></span>.</p>
</td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Ge systemraden tangentbordsfokus. I översiktsvyn <span class="gui">Aktiviteter</span>, växla tangentbordsfokus mellan systemraden, snabbstartspanelen, fönsteröversiktsvyn, programlistan och sökfältet. Använd piltangenterna för att navigera.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;">
<p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Up</kbd></span></span></p>
<p class="p">och</p>
<p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Down</kbd></span></span></p>
</td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-workspaces-switch.html.sv" title="Växla mellan arbetsytor">Växla mellan arbetsytor</a></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F6</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Bläddra genom fönster i samma program. Håll ner <span class="key"><kbd>Alt</kbd></span>-tangenten och tryck på <span class="key"><kbd>F6</kbd></span> tills fönstret du önskar är markerat, släpp sedan <span class="key"><kbd>Alt</kbd></span>. Detta är detsamma som funktionen <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>`</kbd></span></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Esc</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Växla mellan alla öppna fönster på en arbetsyta.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>V</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-notifications.html.sv#notificationlist" title="Aviseringslistan">Öppna aviseringslistan.</a></span> Tryck på <span class="key"><kbd>Esc</kbd></span> för att stänga.</p></td>
</tr>
</table></div>
</div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h2><span class="title">Navigera mellan fönster</span></h2></div>
<div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F4</kbd></span></span></p></td>
<td><p class="p">Stäng det aktuella fönstret.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F5</kbd></span></span> eller <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>↓</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Återställ ett maximerat fönster till dess originalstorlek. Använd <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F10</kbd></span></span> för att maximera. <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F10</kbd></span></span> både maximerar och återställer.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F7</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Flytta det aktuella fönstret. Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F7</kbd></span></span>, använd sedan piltangenterna för att flytta fönstret. Tryck på <span class="key"><kbd>Retur</kbd></span> för att avsluta förflyttningen av fönstret, eller på <span class="key"><kbd>Esc</kbd></span> för att flytta tillbaka det till dess originalposition.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F8</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Ändra storlek på det aktuella fönstret. Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F8</kbd></span></span>, använd sedan piltangenterna för att ändra storlek på fönstret. Tryck på <span class="key"><kbd>Retur</kbd></span> för att sluta ändra storlek på fönstret, eller på <span class="key"><kbd>Esc</kbd></span> för att återställa det till dess originalstorlek.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;">
<p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Up</kbd></span></span></p>
<p class="p">och</p>
<p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>Page Down</kbd></span></span></p>
</td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-workspaces-movewindow.html.sv" title="Flytta ett fönster till en annan arbetsyta">Flytta det aktuella fönstret till en annan arbetsyta</a></span>.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>←</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Flytta aktuellt fönster en skärm åt vänster.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>→</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Flytta aktuellt fönster en skärm åt höger.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F10</kbd></span></span> eller <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>↑</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p"><span class="link"><a href="shell-windows-maximize.html.sv" title="Maximera och avmaximera ett fönster">Maximera</a></span> ett fönster. Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F10</kbd></span></span> eller <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>↓</kbd></span></span> för att återställa ett maximerat fönster till dess originalstorlek.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>H</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Minimera ett fönster.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>←</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Maximera ett fönster vertikalt längs vänstersidan av skärmen. Tryck igen för att återställa fönstret till dess tidigare storlek. Tryck <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>→</kbd></span></span> för att växla sida.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>→</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Maximera ett fönster vertikalt längs högersidan av skärmen. Tryck igen för att återställa fönstret till dess tidigare storlek. Tryck <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>←</kbd></span></span> för att växla sida.</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Blanksteg</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Öppna fönstermenyn, som om du hade högerklickat på namnlisten.</p></td>
</tr>
</table></div>
</div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="a11y.html.sv#mobility" title="Rörelsehinder">Rörelsehinder</a></li>
<li class="links ">
<a href="keyboard.html.sv" title="Tangentbord">Tangentbord</a><span class="desc"> — <span class="link"><a href="keyboard-layouts.html.sv" title="Använd alternativa tangentbordslayouter">Tangentbordslayouter</a></span>, <span class="link"><a href="keyboard-cursor-blink.html.sv" title="Få tangentbordsmarkören att blinka">markörblinkning</a></span>, <span class="link"><a href="a11y.html.sv#mobility" title="Rörelsehinder">tangentbordshjälpmedel</a></span>…</span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-keyboard-shortcuts.html.sv" title="Användbara tangentbordsgenvägar">Användbara tangentbordsgenvägar</a><span class="desc"> — Ta sig runt på skrivbordet med hjälp av tangentbordet.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
