<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Launch a restricted guest session</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="user-accounts.html" title="Användarkonton">Users</a> › <a class="trail" href="user-accounts.html#manage" title="Hantera användarkonton">Accounts</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Desktop</a> › <a class="trail" href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Launch a restricted guest session</span></h1></div>
<div class="region">
<div class="contents"></div>
<div id="restricted" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Temporary session with restricted privileges</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Once in a while a friend, family member, or colleague may want to borrow your computer.
The Ubuntu <span class="app">Guest Session</span> feature provides a convenient way,
with a high level of security, to lend your computer to someone else. A guest session can
be launched either from the login screen or from within a regular session. If you are currently
logged in, click the icon at the far right of the <span class="gui">menu bar</span> and select <span class="gui">Guest Session</span>.
This will lock the screen for your own session and start the guest session.</p>
<p class="p">A guest cannot view the home folders of other users, and by default
any saved data or changed settings will be removed/reset at logout. It means that each
session starts with a fresh environment, unaffected by what previous guests did.</p>
</div></div>
</div></div>
<div id="customize" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Customization</span></h2></div>
<div class="region"><div class="contents"><p class="p">The <span class="link"><a href="https://help.ubuntu.com/community/CustomizeGuestSession" title="https://help.ubuntu.com/community/CustomizeGuestSession">
Customize Guest Session</a></span> online tutorial explains how to customize
the appearance and behavior.</p></div></div>
</div></div>
<div id="disable" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Disabling the feature</span></h2></div>
<div class="region"><div class="contents">
<p class="p">If you prefer to not allow guest access to your computer, you can disable the <span class="app">Guest
Session</span> feature. To do so, press <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>T</kbd></span></span>
to open a terminal window, and then run this command (it's one long command, even if it may be
shown wrapped on the screen - copy and paste to get it right):</p>
<p class="p"><span class="cmd">sudo sh -c 'printf "[SeatDefaults]\nallow-guest=false\n" &gt;/usr/share/lightdm/lightdm.conf.d/50-no-guest.conf'</span></p>
<p class="p">The command creates a small configuration file. To re-enable <span class="app">Guest Session</span>, simply
remove that file:</p>
<p class="p"><span class="cmd">sudo rm /usr/share/lightdm/lightdm.conf.d/50-no-guest.conf</span></p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="user-accounts.html#manage" title="Hantera användarkonton">Hantera användarkonton</a></li>
<li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="user-add.html" title="Add a new user account">Add a new user account</a><span class="desc"> — Add new users so that other people can log in to the computer.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
