�PNG

   IHDR      =   ڲ��   �zTXtRaw profile type exif  xڍQ[!��=>8���Io����I�N�,�Н�����qH9J��`a��A��:�@ 2u�5X~��24�T]co��%~կF+�E�p�(�����b�nd�ϛ�VkDh�x�9���6Z;`G�S��O��)E�8#p�}�n���(���+�W)�'<IH�=�tI��v���be"�O�O�Թ�Ɨ�ڗ���{G?��X�.Tvwd�q�  �iCCPICC profile  x�}�=H�@�_S�"�q�P����U(B�P+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�F�iV�,�鶙N&�lnU�"�D0Qf�1'I)���{�z�Y���}j�b@@$�e�ioOo��}�(+�*�9�I$~�����ό���<q�X,v����dj�S�1U�)_�z�r��Uj�uO��p^_Y�:�a$��%H���2*��U'�B��>�!�/�K!W��B������w�Var�K
'����B�@��8�ǎ�<������W��'���;����붦��;���!��+i
��~Fߔ"�@��[k�@��J� ��h���}����ۿgZ�� ��r�(˞�  \iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:2d9e2d3d-0606-44c7-a2e6-8851d0aae043"
   xmpMM:InstanceID="xmp.iid:8d40663d-d604-4a43-9768-72b9782addb4"
   xmpMM:OriginalDocumentID="xmp.did:372531c2-3675-4fea-b0aa-fc39f464d3ec"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679601280017888"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T20:54:39+01:00"
   xmp:ModifyDate="2023:03:23T20:54:39+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:904ca2ad-0826-4c2c-858b-1328950f0947"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T16:28:11+01:00"/>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:5f8a3a89-89d5-428a-9e61-0f427ab1d562"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T20:54:40+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>+Z �   	pHYs  �  ��+   tIME�
*==   tEXtComment Created with GIMPW�    IDATx��]{�UU��s�s������z�<4"Z���*5R��H31�,M#�ife�F��GJ��G��`Cq��Y��20��T4!.�@���}��k�5���{)�5��.��k}���&@�!B�"D�!B�"D�!B�"D�!B�"D�!B�"D�!B�"D�!B�"�G bKK"�/�q���NN�!B����_��u뺻�_���>��[Æ0`@]��O�>�rȒ%K�(�ӧ��#�������������8�����8 :;;�Ν��٩~w���s�έT*������WÇomm�K�;�B�����k�㎩S�FQ���v��v�ms��=z�84q6����g���2q�ąΟ?���t��WS�L�я~���E�ԩSo��[n�eܸq��?!B��oƀ*�
 ��߿o߾>_ikk����G���������pSS���J�㎻�;�����{�q��͙3�C��Ϡ������L���^{M�4)��<p��v�?0cƌ3�8 6n�x���oܸQ���5k���m۶�{�_|q�Z57q뭷w�q�v	b'�8��:꨿������?f̘��>���ӧR��򗿌�������Z>:bܸq������8bĈ��=�ܳ_�~,�뮻^��j�:r��t��s�=�O�~��V*�j�:~��E����gƌ᪅��Eww��m� `ӦM[�l)�|{{�W\1a8�G�}��n۶mذa�ﾻ�+GqĬY�^z�w�y V�\Y�Tn��=�أts�c;v�֭[�̙3a[o�����J_?��S�?��r�!|�-[~�ӟ�y�/�����iӦ�^���o~��G���/<��sG}���7o�|�%��x�'�pB�>}n�ᆖ���#G�w�y ����~��&LX�n�̙3���.�����oܸ�.�S���x��w����[���&L<x��/�x�5�tvv: ����������c����w�y��g�=�cV�\9cƌ1cƜv�i��������ΩS�z����{�G~��Z�jՅ^���>e�]v�����f͚�+W�]�v����;w�I'�������_��s�=7~�x زe˅^�y��_~�;��N[[ۚ5kbǊ�o�}��շ�v�!���o8>��.�̜9���x���g�}�O�~�Yg�^����k�ʕ��9�ŋϜ9����^�r�7���{���O���ܻW�`�q|��/_���{��o���� :;;�;％>��c˖-{����J�2t�з�zkÆ�~xgg�!C֮];dȐW^ye����>��m�����~饗>��#K�.=��s_xᅕ+WΟ?�����G>r�i�]u�U�J�SNiii9��#�,Yr�=���)D�%�l�BD#F�0`���?OD��3g����-Z���o�8p������Q�F�3f��ٟ�ԧƌ�|��o��[n�6m�^{����:f̘�~��'�T��bŊŋo޼9e�ƍ�8cƌ{�����+.���U�Vp�C�y��G�On޼�R��;�����U��%bG��N;m��ٳgϾ��+�N�
 �^z��^���.�L��SN2dH�C��o�뮻�9r��������.\�y��e˖�~�� �z�꧞zjܸq��Y���ڎ=��c�=v޼y�0a  �W��7�|���߰a�ƍ׮]�R���.<�#&O���㏯_� 6mڴ~��u�ֽ��Ç�����g>3jԨ�^z������^�j�o�1bĈA��s�9�Je͚5Q���;�g�^�xq��B�؁b�}���ˮ����~�W�?��SO=���.=zt���˗?��CK�,Y�l��?�lٲ�������O?���D[[[Z"��/�y睯��{�?��'O�<q��+V|�s�#" 4h�����+V�;�����c�immEĉ'�|�ɳf�ڴiS�^!B�@�|��N ��k�Ν;7娦N�گ_?�!�t�p&�c X�n�c�=���ڬ�FKK�7��6L�4�裏�������җ�4eʔ�o�y�֭TKy䑳�>{���3g���[�nmkkkmm}����~��s�>��S���ƍ�nݺ�n�577�X�b�֭����6mڴiӦQ�F�;)D�q�����/����ׯ_�$Ç_�nݪU���j:`��555�|��k֬����'N���*�������8����ׯ_?bĈ�7�����������k��f͚u�����/8p�A�ZZZF���_�jܸq�\r�����k�555�8B��^�x`�]w6l�����5k�l۶�o߾p��)Sn��^x�������뮣�>���#%��<��6��������ݶm��w�;��|���)���<�����^8��/�|Μ9��� p�QG-^�x���{�g>��OO�6m�ҥ���I'��dɒ���{��k��6d� �?��E����7~��+V ����s�]u�U---ӧO��o~s�}�]t�E 0mڴŋ�q����~��O�{ｓ&Mʿ"D�(n����_�-z�駿�����~O>������K�~�[��	�k����+�lnn�3g��_ =��Yg�u��g/Y�d�����ǌs���ϛ7�����������������|��J�r�UW��X�t�T�VG��'Ǝ���O�%�˖-{�7�y�'�x�c�X�d!B�(q�Wtwwwww�Z�j��� p�	'������o��f�l����~�7vww��=��>��O���o��ɹ�Ɍ	&����5kVJ6z����{��5��c��vkooO	������������Ζ���}�vuu���T����΁V�աC��e�He�MMM)��x�=��}��S'���������6 hnn<xp���g;;;���7D�;P���òhooO]Z���٩VD0`���8p��t(����߿sssWWWGGGGGGSSSkk�A�̭455uuu�[2d"���vuuuuu���_�|gggE 0L�`�"��g���"�FS�N�_IUY�hkk{��r���M�����_�����ӟ��dɒx�4�"D�!B�0q�嗧X��W_M��ɓ'�]����{�ڵ�&Mr}�����vuuM�8���G�뮻�K"D�!B�"D�!B�"D�!B�"D�!B�"D�!B�"D�!v��~�_�^�����W �jP�o�>� X��oQ�@X�.*�C@ ��`�߼�1�@�7���l7H�+݈5� ����D @GQK�Z�Z&�_#�����+GK�"~�ҏ#QzB )v9;��L��D���p1�o L��� (! �����D���b!ж$I�ԓ�Rv*I�GE��j_Q�bzhX��|[�=�~��*�?�X�9T ��a����;�]��?P9����oH��I��@sC�V�_PN����1,�d�D����pq@�w�=W��s"�$��]s����V����W��m�t���|�aG�C~Ay����������3�ϝzf��g��H�y��w	�Iȏ-���wP?W�1��~J�o[��&姊QC���'2�*�
���Ko޲d�Q���r����ɨ�?�M�+(\H}\ �F#�4�c�:h����wɿ#�]X��а�j5U���A=�&�T����1(>L��I�L
��s�OV��t�A@ 	I�8{��H�X��X�=Ǩ���]�2ˊ[F�J �]]��C�������
��C���..Q�M�1J��
�����҃j]i�K��{�j/���d���+�8�![	�!��?��/9wT��-��u���KX��r9��J~��cH�|��q�E8���DN<]7�v���u@W;�B-�D�EBT��R2�$A�2��ȉ�Fs;Hh�q�Wk�3�V��"�(1 ���`�}e{���x��Qc���;X�ǈ@D����B"��F�h��~� y�V����˘hܵ���QAW$�]�����M�U�S5�Ő�~�`�]�i�%!�|9�Ъ8"�0���m�u֪ʪt���6���e,7=���1I$������-GM��Fַ�XN������ߕI �4r]�W���I�B�u�V��(S	6��s�E7���d��K�2�)�m	T"�D���^q,��qSq�����Q�O�����T����	�2~%`@�"e9Am�F��I�8�oɧ(M[b1a��(�%>�PN%=�aȒ��Y"S]�gd�>�?��d_�J���T���h�R�TL���$~R��ŭ����B�8��H��>iA+ۄ:�`c����h叫�xE��O{6�)�Fb�.�V�!/ �;�����̃�t�Y2�iA�P�$�o���5�<*��Lt�+r5��`�j@�@K��n2�GQ��T�|w6��j��C���K$�0�AT<�$ɪl�U*�Ja�ҩ���@���}Q����OZ�Yư�[	Q�.-2� ۘ���4����9�#rW���B1?�XЌ�-�%]��yVѕ
�
p@�+��t��O�wZ�F\qT�W�J&��wu`�$BX7�Rpz�l��r�N�a�牿톰$���+��'�@A�P����$߫.�����ҙ=I�hu�w��P|�����eIFNqB�E"�7eŅ2T2:E�M�j#��@�\\OqU#�	���(�H������F�M�*�Rs��b��,���� ])w�]�s�&C6�M�d�+����"��ntvt�^ �Bu�ϕ��҂P��\�e�?��an�:6�T?��\������8�Ľ�=�Yt�^���"	�U}E~�����)$��1�䠈��x$�ߐ��N2SP�M M�&���w�`��b�ҫ;
�"�ՠ�c[q��般�˅�W�w`s\�`�~���۬$SE�~��o5wC%��Ф���"�O��+"d��`a�X�a���4$!%=�����E_��+4�Iܕ���@��fъi�t�9�r���!x�+�]���S�W��+��ˠ����
]'����&�G,���b�ቚȲ��/j��E�D�����*�׶�T��m�ZR����U9��ћ�ۈAP&���Й�~y��Ucsq�� �ey��l� ��"@���F�R=�l��1j�+1���2��T�:���*��f� q�D `�V�x�{��%**��T���.�"O�v~�Dd�+�r� J�
�q��^ h�JЕ�!GZ��ЕL\AI�`ω+����ZA�Ъw��hV�I�a�d���?���r�K���W�f0�cӶ���� +y5S��)�/]��epC��}�C$Y=׹Fk�)[;�E%�(ٟ)�'1
���GS���P~�&%yC�Õ(j�*J5��vK�Oā#?�V�\{��M�y��,�@+W)��8o�4m���u�V$mE�a�"��.mM��BW���6^A3�"�ze�"l&&���tt���E=��5�3��CW�+h��^��׋!ӳS	�2��
���v~4�P��Ъ>\��3ٙ 4�,�S	��������R���4}%N%�J���ꈖշP�`'��s��^���F�ƒ�]��,'T�-X �9I"�=���KQ��T��o\����+�*힥�SH�OY�!�B%m�����"�Tu�0��*CMaV�RI��d$���j�͆�����eCW�c\=���ȧ`�t�ٕ�ut��.U(t����Ć�21�H\��ŀȊ7=�+�2�k��z�)g�L6����m��ՠ�3��$�歨��@^���W�B��S�v�ʴm�rЁ�먼�FW���\�vv�o� �kM�M���2T�/����,O����qS�h J:�,@�B�n��M'�J��s��Xa��"�j�D[�
ާl�-Xf�OD�<����l��д�+��
e~&?t���Rt.t��h}��ӥ�uIک��B���~t%���
EE�!��zW��w�a��a����J��E=�+�N��8�m{��V9�iڮ�A.����׫N�P��l���S^J���1��tߨ˗�<p�+)�+�(���hR`���zM�Nf��_j6T�k:��(��Q(5"�^�b6M'��z�#+G*�`�,�d݊�؉`c�A��+3:��+�])g�С�����^BW�.���(u��ϋ�!��z���s�vh%��R\�%�*�5CX�j�B���n���F�y�f{�m'>��T�-9h_��Ӵ��Я���r�Q�������J�X�O��S3�T�G@��"�BN��T��q�%�H�+�h�:�B:���D"M	�P>��Bh�Ϳx�A�!����f�z�C��{����6�s�@���P���,�+(官�T��Q?[��aS)*S�:�+�DO�9Еӥ]Nj��N��t� ��M\9��b��|��i	��u^dU�;��mf���ӻI&ɝ�G}>|x�W�C��s�{��7mw���A�A	��f�+9��;��������B�q*l�ey��_�r�6]/O�c�\��j����*��.��-;�I1���2s���T�L��$.!�����gMb�d��"�ڀ��D�3'y��Z�����Gn�`�+H�Dcō�Ҳ���]�0{���mTy/�Q���.�+��2|D-
'�8:@��|^�X�LqUJ\i>�V�\�%���w-oA�Q�H]��*9.����Wnk�2|�-\[Q�y��qO�xh��×�>+�SՋ�W]� �e���:��Y�i����;��C�^�K'Bl�T*�<� �Pa���<�.�0�Ic���^͢�����*)�'��g�;��=d�5?dCiA>j9�8@S�Dr�RB��Ay�2���	+Q)-�c��D����C����̑K��EYU[ѕ��z1�]t��@�׈�h%�YHt�p�3ߐ̾�0-��Z��n��gSfA�G�8�2K]�oSg�d�Sb+*���ea��ѹ��
��Az���W\�_t;r��1��s��A�|q7�qպ�F�uϷ���	������FDl	9�CM���B���d愢9��OI%挨tXt �\���x{��RE�cR�!�1�2.c>�8Еv'��ʄ9��DW���*�ӊ��L�Ns2L�K�l/���B�E�r+���|UCXhCZd\�lzZ�Wjnbs^p<��CsDm��2G�Rm��+X�%��o�i;Z���WrK�2wGr��ȥ^l8��;��vXэ�th �WC� D���~�M_��(��b�f^�E�A���Jv"9=������B/;��幡�T�b�Kk�E�-��e���]d]�II��Z Z�5
�E����j���2GCW�m�]��+)���2���
��J쁣b��CW6;xT~�JR	q���F\Y����v�X`�8�a�Z�4���z=[rQRhu΢$ҟ|y&-��#2�
s7�6�`�^9��䩧��PzePgN���1,v&�͉v~�;E&T��(�����铺N�j5�d3����,R8�eB�����5���b#.�.O@�U7Q2��@�.T�F!��Z�hc�:ځ����*>3P�� ��G�Zj�4t�
���B]q�R��Y���r;rE��ǳT{ˁ�zC��"�L1�ON����ł�T�T�e:�E@�[���4��tG��mwY3���"�(�4�%9H�@�X|H%�z.�*EH�Cz2�;	�U� ��E��LְW.yM�	A�*bu�M  U����[�S>��@�Mų��JZ��ms�)�ku�Ū��	԰�_�%G�4�v򑐲�EJ�/�.Ec�F$�,zͽFsHj?�]��t]	�H�����]���$Ā ����Q;�^&�+՜LFW=�c��jA�Ƃ��.U\�9���h��?�D^����^����D��V�
˶/7uvڊʕ���sP^���^���WmWO��P�t��H&�2�j jϸ�yU�Ί���K���fJҬ)����U�4  IDATMY�oMr+��9������
��m�4�z��	�j�e4�$�(G��RcGR�>_]��MIŚ>�G"�ӈ
,��CZ6P�5?O?I�k����\�M��� ��]�.��W���L�%�+��`DtU��.���CWZ�Qj,(���=A�;'h�V(�X�Yl���Ĩ�N��~(���w�i.Z�BX��fKH�ي��ˎ���/C]pʁ�n8h��]Q����ZW�ꓞ@k��zb.p�������B��8�DQ��T�:�'���ـ�ͯ(_��}���Bs �%e���i)N�Q'.�B4(D$������#N=����&pC��*�X�)Kt�̧��(�\b��2�v����D9|�ƚދ�7��(�ѕ\>����k$�1��+^Y��r�i�zWn%{	���(�ނ�%]�ݤ:���J)���Ȣm�k;h.AŮ8>�����4�3?l�ep؁�=��FW_��tUW���)��,�$�I[Fh�*�e���R?�*��3(:����?��m�&�+QT����8Qq���A� ��=��Ш�&L�Y�x&�7�'V��Ptq5 ,1F�@urj4kz����*�a��;��@^U@��@$�Q$|ɜ��%1����ȩj'˰����PnJh7jg`����fW��J��b3k�D1��,D��8�X+�*����r�հh���!�#U��`]?Z��ͺ9������VT��d�^�����2@C�Ai>��-��`�휩���z�w`�􆑉+]��ّ�O��Fb��M���J���
�O�}���Roe���H�6a�T�c�J��lX}��Xd��N� �e�2�c��T�V�M(���FMWշPHm6Ӥȡ���\����^_�,]�����-�MmfW�6�(�1��@��w�7Е�`�Aѕ��r����+1'h�V��,ڃܠ�*l<���t$A`�����p�W�������ʠ�\����Ŕ^�[zU�/ٰ��v_V�����}�XTvo����=�ʓ�dO�FR��y��=
ĈMq���I���������|\HN��<o�!��r+�bMq� >�HY���� �'��o�0I-�I9)��(�8�F���	5���5���.�[�}��P5mp@FWH�<
�խi���?J܀���qFoK�Ut��#�Ջ4@�iA��'ffi`���ܸ
{���2����K+�p�,�K��W>�A>�c�M��1���6Ѵ]�J|�W�^"Zp���돈�;����<E��� ������"5'`cm���r�Qs\)z �&�Hr�#GQ��y>���G �%a�|�P;��4;Q�����	�	�@�1�J���P�8DҒ4�7��xP $tŪ�P/:d�gjSq��
YoJ4��G�Qm�G¾��(2�򉖛]��
et�5z2ѕ�L��+O�U^(��ƈ+����r�*qq!�W���v�=����8+�z��"s���m��$��!�R9(��Eg���Ђ?@(�VЕ�m���zEVB��S�LH�� ˵sv�ѕ6\8*������qتFqS\�����.�2#I荈H�u�ޡ�%Y�#P�3�����K��R7d�[4 
��|6Jḑ&Ӑe[)���9�q3�(k�&��WD�i��X�8mp�Ր��Q0�U�|����3��0�H2iD�ev���qu��+�v2l���O�NW%Ղ�WV����C+WQ9��	�k��R#^��'E`1��-��E	��� ���[�����������6�z%�+({WsF/s,��t�3 ,�s�<�/u�X�+y9#�ɺi�1��q5�te���N@B�c���B,�_"qqB��J�hP�N���^,n匨!SoQ�ֱ&�/p!gD�����P7) ����F�����9��z�}x0���;[�*|��b2}*B�ʝ��֡%(�(��z��LBN��BY!�Oai�R#�����rB+1�\Z��f���^��k<�m�d*���N[�M;u*%�˴�T�y���tn�vp$���ė�ǮW����h��S4���`յ4��̌��XB&H��-��mD�jU���5h,��\��tL��&�P�b��\@c�<�����F1K*"sm$���X��� Q�%�BK	�|4ML���T�p�%�@��Hd��[&�Ux�A�ȠZ�h���Y���">��a=we)d0Bsɗ���7��Pt��F���b����y)�ʈ+Z�I�Rr��E5���a=�[�^�"������"�׶�m|E��Ѵ]�~�ut��28�W<9(5t�_�q{�I����ݲ��3 ,��LҘ��Dԟy�?̙eCdu�A�>q\��枥�5�����7&�}"�B-)��B5�}�K�Pn�1i�Ʉ�?8�*\݊��f�9V�*fЊ��v����-4���Z9��t��x��޲�OJXN��v=�s ��&��b���D**0�̥���"-��v�	]e\��6-fW=GW�^�y���J,t:��`���<��0���Aem��#bSb�u #���#Hu�&\�����W�%9�0m���5_Ғ�?�eԗ㚔���������;��c���:�,�$�ȇ!"iQI�Wb�գ��:���Nͻ�?' B�E�h��W�>Z�h�ذ�C2w���0&�Gf��� m�ѹxʕRXC
I���U
Rq&�M�KE�j*�H���T[^L��Y��V`s��7��Y�PF��"�
"�H2\ "{d:�ѕe�hCW��;#�7;j��j��z%�&�2qB� ��Z�B=;��U��Ї��+N�X+�O��PM5H_Y��fa���]����|��jX/�����}O���������;�v��3�z2XGl�VZm�[zhZrf�ܵ#��*��m6Q� c�����j�PM���"BA|�J� �����B\�?�SAj�?$y�$�a��Ј��u:�v��#Qq�P�d*5ۇ���M��C�,KQ����	Yfs��&
ɼ�TZ��9�)�v�ѕ
��H��}�t�+�4�ǔ�����k�
$�~��|��＞,M
,x#����$���Gld"k���M_�8/�V������p8�	X���FW��y�.a�_K�S�79h�s�r��<n>�pZ�Ja,٩,�NL��� ��W�-�[�2A���+�S�M���O��]��9kMC�"G����"y.�N���?H�Ƥ@�QF��\�����cD$�c�v�
�F�=�o��֎I�B�H��k|��">�F�ۀT�B̻!�p%���@��t,��]���PN�eIGW�F��>�e�^/�hzva�����VE����x_�'N��(�X��%��N���l ��b#������<9hdZ�SLΌ���EG�'��k8��y����%�{��)0����2 o(�@+�����9��֕(�W��K��meN�P�[�4C`XJ�F����F�sx�	���̄�0�qX&�i��SKҴ ��D1��Hj��E���gy���*� !R^'H	08��#R��`*%����AM��ܠ�+U�m����i���@W��
�uiG���^��T=;J���+,9�����t[��(k1A�T��F�+���6Z���~�%�C�|�_wK[�ANҚ�C��A�:��=�CC�j�����3X�+*�*q�7����H��J\CW�	p��F2�1�������T��S��)��'<�YԚ-�pqgPN�掖2=H��w1���a�2_*T�@�p*EW	0���_b32��^t���,EW��^SMC�:�j&�J�lD��IP�v&�Rd�)�<F�`*�l��wɎ� Mҥ���д����J����tO//�R#���gX�d"�*�S:0��0YH,t�τ�գW p����ʬt%��;p�e+�h��AYz��+���\���d��^Y�9��%te����;�%�Q��?CBn�i�8R�>Z��jTa�<}#ʈ��+�t���Q����R��U��<��̛73tE9�B�3�[�|1ŕHx%f6��O�r�Y	"�> �D� ����L�p't�i���d%���y5�QD�O=eZu$ҐD�(b.��)$Ս��Ħs��H,� ;@g^�+	[����� ƹͮ�v����� �+S0f5E�!�����Z�����Ppv���J��<�W��V����*�Lۥ]%����+�^��z��8f5"GW���f]�T(|�,�4�-��L7�2	b|o��G�nř��ڳ����FBeb�_��@���5��[F��sR�nd$�a�Μ�fd�V
l��51_{%���x��9/�$����O�R��,�K�YR� $��O_�h����Hi�������9�0���!���T�O�4�����M(l=����68�]�@�bGW���D�y,uW�-*�VXNZ�c�g�Y'y@��W{B2}U�vЖ�rkx�>�����[�=9ؓ���sVA<�:w.t~�����b�`�ʮ82�X�b���'.t!T�8���������Iԟg�W��;�gLQ D�N
��{"��4�Ө�����#s�P�k�""��Nꠕn4)���S�8`�֊��!l�&� �*
d`�C�K��EPK��R�E{�Z�V\��N�P�� ��ЕD�� �I\�E�J4߄]�EW�*�K����P"��ѳcA7�B+�zC���@���� ,qg�f�N���-9X�E$��ė�H��2�/���'�x��z%��͛�\-��w���u{x����!���U�q�.���r�u"���#�W����v����S�؎�Բ�X=f��m���W�CIj:�g&i����H2e��3����j�iG�2e1���D0��y�MC
F�?B����H�V�ȮV~7�����G1'�2S3D���R�Z��A�|��!7R���H!�$�T��~u�+���IڡLtE����]4O7/xd�Z�\�&���Ba�ۖ<�7H_�{R���'�-z��}:j����F�2�̳�Kz%�[wOQ/�b�XHX��	Rg���U��*+��@A�#nJPh;�>���4A��CYa� � 1�	ҏ�4�J�g��+���4GR�_V~X�T����9@�$��<B3>��A���*�*q�H)T�1b��9PJO?qvQ�G���b�E�6U#W�
��-4�i���ق��!��52�V�HRV�AQd�mP"��նٖ��	
��AYe�z��C݇��5�D �>N���:Y��]߀=9hEW���Ά~-q,�Sl�C>�+39艮z�STDWT7��Rt���S��y�fI揄K�1D}�8R[�	1R4C*9�2	�~���[;�~�n16[ ���Ifu��<�#-�u�A&�"��)$��Q�V����ۖ���W��V�nf�3�X��<7�P�.4�R�xa������IH��⇈㰢a��E�0�Hk��_�\����� NlI���*�R�Dy��l%j��+h]ټ�l���'-�wC+4AU��N��F�}�ޠ�uJ�+���������V9�H)X*-���-q���i�˰oҫ���W�.J���
���y���ާ��.9z0i�;�    IEND�B`�