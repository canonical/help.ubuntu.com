<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vad betyder ikonerna i systemraden?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html.sv" title="Ditt skrivbord">Skrivbord</a> › <a class="trail" href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Vad betyder ikonerna i systemraden?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Detta avsnitt förklarar innebörden av ikonerna som finns i det övre högra hörnet av skärmen. Mer specifikt, de olika varianterna av ikoner som erbjuds av GNOME:s gränssnitt förklaras.</p>
<div class="media media-image floatend"><div class="inner"><img src="figures/top-bar-icons.png" class="media media-block" alt="GNOME-skalets systemrad"></div></div>
<div role="navigation" class="links sectionlinks"><div class="inner"><div class="region"><ul>
<li class="links "><a href="status-icons.html.sv#universalicons" title="Ikoner för hjälpmedelsmenyn">Ikoner för hjälpmedelsmenyn</a></li>
<li class="links "><a href="status-icons.html.sv#audioicons" title="Volymkontrollikoner">Volymkontrollikoner</a></li>
<li class="links "><a href="status-icons.html.sv#bluetoothicons" title="Bluetooth-hanterarikoner">Bluetooth-hanterarikoner</a></li>
<li class="links "><a href="status-icons.html.sv#networkicons" title="Ikoner för nätverkshanteraren">Ikoner för nätverkshanteraren</a></li>
<li class="links "><a href="status-icons.html.sv#batteryicons" title="Strömhanteringsikoner">Strömhanteringsikoner</a></li>
</ul></div></div></div>
</div>
<div id="universalicons" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ikoner för hjälpmedelsmenyn</span></h2></div>
<div class="region"><div class="contents"><div class="table"><div class="inner"><div class="region"><table class="table"><tr>
<td><div class="media media-image"><div class="inner"><img src="figures/preferences-desktop-accessibility-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Leder till en meny som slår på hjälpmedelsinställningar.</p></td>
</tr></table></div></div></div></div></div>
</div></div>
<div id="audioicons" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Volymkontrollikoner</span></h2></div>
<div class="region"><div class="contents"><div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/audio-volume-high-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Volymen är högt inställd.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/audio-volume-medium-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Volymen är normalt inställd.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/audio-volume-low-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Volymen är lågt inställd.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/audio-volume-muted-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Volymen är tyst.</p></td>
</tr>
</table></div></div></div></div></div>
</div></div>
<div id="bluetoothicons" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Bluetooth-hanterarikoner</span></h2></div>
<div class="region"><div class="contents"><div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/bluetooth-active-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Bluetooth har aktiverats.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/bluetooth-disabled-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Bluetooth har inaktiverats.</p></td>
</tr>
</table></div></div></div></div></div>
</div></div>
<div id="networkicons" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ikoner för nätverkshanteraren</span></h2></div>
<div class="region"><div class="contents">
<p class="p"></p>
<p class="p"><span class="app">Mobilanslutning</span></p>
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-3g-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett 3G-nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-4g-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett 4G-nätverk.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-edge-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett EDGE-nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-gprs-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett GPRS-nätverk.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-umts-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett UMTS-nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-connected-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett cellulärt nätverk.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-acquiring-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Erhåller en cellulär nätverksanslutning.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-signal-excellent-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Väldigt hög signalstyrka.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-signal-good-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Hög signalstyrka.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-signal-ok-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Normal signalstyrka.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-signal-weak-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Låg signalstyrka.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-cellular-signal-none-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Extremt låg signalstyrka.</p></td>
</tr>
</table></div></div></div>
<p class="p"><span class="app">LAN-anslutning (Local Area Network)</span></p>
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-error-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Det har blivit fel vid sökning efter nätverket.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-idle-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Nätverket är inaktivt.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-no-route-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Det finns ingen dirigering för detta nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-offline-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Nätverket är frånkopplat.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-receive-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Nätverket tar emot data.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-transmit-receive-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Nätverket sänder och tar emot data.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-transmit-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Nätverket sänder data.</p></td>
</tr>
</table></div></div></div>
<p class="p"><span class="app">VPN-anslutning (Virtual Private Network)</span></p>
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-vpn-acquiring-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Erhåller en nätverksanslutning.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-vpn-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådlöst nätverk.</p></td>
</tr>
</table></div></div></div>
<p class="p"><span class="app">Trådbunden anslutning</span></p>
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-wired-acquiring-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Erhåller en nätverksanslutning.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-wired-disconnected-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ej ansluten till nätverket.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-wired-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådbundet nätverk.</p></td>
</tr>
</table></div></div></div>
<p class="p"><span class="app">Trådlös anslutning</span></p>
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-acquiring-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Erhåller en trådlös anslutning.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-encrypted-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Det trådlösa nätverket är krypterat.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-connected-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådlöst nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-signal-excellent-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Väldigt hög signalstyrka.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-signal-good-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Hög signalstyrka.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-signal-ok-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Normal signalstyrka.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-signal-weak-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Låg signalstyrka.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/network-wireless-signal-none-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Väldigt låg signalstyrka.</p></td>
</tr>
</table></div></div></div>
</div></div>
</div></div>
<div id="batteryicons" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Strömhanteringsikoner</span></h2></div>
<div class="region"><div class="contents"><div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/battery-full-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är fullt.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/battery-good-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är delvis urladdat.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/battery-low-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är lågt.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/battery-caution-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Varning: batteriet är väldigt lågt.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/battery-empty-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är extremt lågt.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/battery-missing-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet har blivit frånkopplat.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/battery-full-charged-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är fulladdat.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/battery-full-charging-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är fullt och laddat.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/battery-good-charging-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är delvis fullt och laddar.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/battery-low-charging-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är lågt och laddar.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/battery-caution-charging-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är väldigt lågt och laddar.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/battery-empty-charging-symbolic.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är tomt och laddar.</p></td>
</tr>
</table></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p>You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
