<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Dölj en fil</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html.sv" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html.sv#faq" title="Tips och frågor">Tips och frågor</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Dölj en fil</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Filhanteraren <span class="app">Filer</span> ger dig möjligheten att dölja och visa filer efter dina önskemål. När en fil är dold syns den inte i filhanteraren men den finns fortfarande i mappen.</p>
<p class="p">För att dölja en fil <span class="link"><a href="files-rename.html.sv" title="Byt namn på en fil eller mapp">byt namn på den</a></span> med en <span class="file">.</span> i början på dess namn. För att till exempel dölja en fil med namnet <span class="file">example.txt</span> ska du byta namn på den till <span class="file">.example.txt</span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan dölja mappar på samma sätt som du kan dölja filer. Dölj en mapp genom att placera en <span class="file">.</span> i början på mappens namn.</p></div></div></div></div>
</div>
<div id="show-hidden" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Visa alla dolda filer</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Om du vill se alla dolda filer i en mapp, gå till den mappen och klicka antingen på visningsalternativknappen i verktygsfältet och välj <span class="gui">Visa dolda filer</span> eller tryck på <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>H</kbd></span></span>. Du kommer att se alla dolda filer tillsammans med filer som inte är dolda.</p>
<p class="p">För att dölja dessa filer igen, klicka antingen på visningsalternativknappen i verktygsfältet och välj <span class="gui">Visa dolda filer</span> eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>H</kbd></span></span> igen.</p>
</div></div>
</div></div>
<div id="unhide" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Synliggör en fil</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att göra en fil synlig, gå till mappen som innehåller den dolda filen och klicka på knappen visningsalternativ i verktygsfältet och välj <span class="gui">Visa dolda filer</span>. Leta sedan upp den dolda filen och byt namn på den så att den inte har en <span class="file">.</span> i början på sitt namn. För att till exempel synliggöra en fil med namnet <span class="file">.example.txt</span> ska du byta namn på den till <span class="file">example.txt</span>.</p>
<p class="p">När du har bytt namn på filen så kan du antingen klicka på knappen för visningsalternativ i verktygsfältet och välja <span class="gui">Visa dolda filer</span> eller trycka på <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>H</kbd></span></span> för att åter dölja andra dolda filer.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Som standard ser du bara dolda filer i filhanteraren tills du stänger filhanteraren. För att ändra den inställningen så att filhanteraren alltid visar dolda filer, se <span class="link"><a href="nautilus-views.html.sv" title="Visningsinställningar i Filer">Visningsinställningar i <span class="app">Filer</span></a></span>.</p></div></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">De flesta dolda filer kommer att ha en <span class="file">.</span> i början på sina namn, men andra kan ha en <span class="file">~</span> i slutet på namnet istället. Dessa filer är säkerhetskopierade filer. Se <span class="link"><a href="files-tilde.html.sv" title="Vad är en fil med en ~ i slutet på namnet?">Vad är en fil med en <span class="file">~</span> i slutet på namnet?</a></span> för vidare information.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="files.html.sv#faq" title="Tips och frågor">Tips och frågor</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-tilde.html.sv" title="Vad är en fil med en ~ i slutet på namnet?">Vad är en fil med en <span class="file">~</span> i slutet på namnet?</a><span class="desc"> — Detta är säkerhetskopior. De är dolda som standard.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
