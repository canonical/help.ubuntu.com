<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använd alternativa inmatningskällor</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="keyboard.html" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="keyboard.html" title="Tangentbord">Tangentbord</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="prefs-language.html" title="Region &amp; språk">Region &amp; språk</a> › <a class="trail" href="prefs-language.html#textentry" title="Textinmatning">Textinmatning</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Använd alternativa inmatningskällor</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Tangentbord finns i hundratals olika layouter för olika språk. Även för ett och samma språk finns det ofta flera tangentbordslayouter, som Dvorak-layout för svenska. Du kan få ditt tangentbord att bete sig som ett tangentbord med en annan layout, oavsett vilka bokstäver och symboler som finns tryckta på tangenterna. Använd det här om du ofta behöver växla mellan flera språk.</p>
<p class="p">Vissa språk, som kinesiska och koreanska, kräver en mer komplicerad inmatningsmetod en bara enkel tangent-till-teckenmappning. Därför möjliggör vissa av inmatningskällorna att du kan välja en sådan metod. Mer om det i avsnittet om <span class="link"><a href="#complex" title="Avancerade inmatningsmetoder">Komplicerade inmatningsmetoder</a></span>.</p>
</div>
<div id="add" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Lägg till inmatningskällor</span></h2></div>
<div class="region"><div class="contents">
<div class="note note-sidebar" title="Sidopanel"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan förhandsgranska en bild av layouterna genom att välja någon i listan och klicka på <span class="gui"><span class="media"><span class="media media-image"><img src="figures/input-keyboard-symbolic.svg" height="16" width="16" class="media media-inline" alt="förhandsgranska"></span></span></span>.</p></div></div></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ikonen längst till höger i menyraden och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">I avsnittet Personligt, klicka på <span class="gui">Textinmatning</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">+</span>-knappen, välj en inmatningskälla, och klicka på <span class="gui">Lägg till</span>.</p></li>
</ol></div></div></div>
<p class="p">Den förvalda inmatningskällan är den som visas överst i listan. Använd knapparna <span class="gui">↑</span> och <span class="gui">↓</span> för att flytta källorna uppåt och neråt i listan.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du väljer en källa med en inmatningsmetod kan du klicka på <span class="gui"><span class="media"><span class="media media-image"><img src="figures/input-preferences.png" height="18" width="18" class="media media-inline" alt="inställningar"></span></span></span> för att komma åt den metodens inställningsdialogruta, om det finns en.</p></div></div></div></div>
</div></div>
</div></div>
<div id="indicator" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Indikator för inmatningskälla</span></h2></div>
<div class="region"><div class="contents"><p class="p">Du kan snabbt växla mellan valda källor med indikatorn för inmatningskällor i menyraden. Menyn kommer visa en kort identifierare för den aktuella källa, till exempel <span class="gui">Sv</span> för svensk layout, eller en symbol om du använder en källa som använder en speciell inmatningsmetod, t.ex. Kinesiska (Chewing). Klicka på indikatorn för inmatningskälla och välj källan du vill använda från menyn.</p></div></div>
</div></div>
<div id="shortcuts" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Snabbtangenter</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan också använda snabbtangenter för att snabbt växla mellan dina inmatningskällor.  Den förinställda tangentkombinationen för att växla till nästa källa är <span class="keyseq"><span class="key"><a href="windows-key.html" title='Vad är "Superknappen"?'><kbd>Super</kbd></a></span>+<span class="key"><kbd>Blanksteg</kbd></span></span>, men du kan ändra den:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på ikonen längst till höger i menyraden och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">I avsnittet Personligt, klicka på <span class="gui">Textinmatning</span>.</p></li>
<li class="steps"><p class="p">Klicka på nuvarande snabbtangentdefinitionen nedanför etiketten <span class="gui">Växla till nästa källa med</span>.</p></li>
<li class="steps"><p class="p">När snabbkommandots definition har ändrats till <span class="gui">Ny accelerator...</span>, tryck ner tangenterna du vill använda som det nya snabbkommandot.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="windows" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ange inmatningskälla för alla fönster, eller individuellt för varje fönster</span></h2></div>
<div class="region"><div class="contents">
<p class="p">När du använder flera källor kan du välja att alla fönster ska använda samma källa, eller använda olika källor för varje fönster. Att använda olika källor för olika fönster är bra om du till exempel skriver en artikel i ett annat språk i en ordbehandlare. Ditt val av inmatningskälla kommer lagras för varje fönster medan du arbetar.</p>
<p class="p">Som standard kommer nya fönster använda den förvalda inmatningskällan. Du kan välja att de istället ska använda källan för fönstret du använde senast.</p>
</div></div>
</div></div>
<div id="complex" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Avancerade inmatningsmetoder</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Rekommenderade ramverk för inmatningsmetoder är <span class="em">IBus</span> och <span class="em">Fcitx</span>. Den senare är standardramverket i Ubuntu för kinesiska, japanska, koreanska och vietnamesiska.</p>
<p class="p">Inmatningsmetoder är bara tillgängliga tillval bland inmatningskällorna om motorn för respektive inmatningsmetod (IM) är installerad. När du installerar ett språk, installeras en lämplig IM-motor automatiskt om tillämpligt.</p>
<p class="p">För att exempelvis förbereda för att skriva koreanska (Hangul) på ett engelskt system, följ de här stegen:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p"><span class="link"><a href="prefs-language-install.html" title="Installera språk">Installera</a></span> koreanska. Ett av de installerade paketen är <span class="em">fcitx-hangul</span>, IM-motorn Hangul för Fcitx.</p></li>
<li class="steps"><p class="p">Stäng <span class="gui">Språkstöd</span> och öppna det igen.</p></li>
<li class="steps"><p class="p">Välj <span class="em">fcitx</span> som <span class="gui">Inmatningsmetod för tangentbord</span>.</p></li>
<li class="steps"><p class="p">Logga ut och logga in igen.</p></li>
<li class="steps"><p class="p">Klicka på ikonen längst till höger i menyraden och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">I avsnittet Personligt, klicka på <span class="gui">Textinmatning</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">+</span>-knappen, välj <span class="em">Hangul (Fcitx)</span>, och klicka på <span class="gui">Lägg till</span>.</p></li>
</ol></div></div></div>
<p class="p">Detta gör <span class="em">Hangul</span> tillgänglig i Fcitx-indikatorn för inmatningskällor i menyraden. (Utformningen skiljer sig från motsvarande IBus-indikator.)</p>
<p class="p">Om du föredrar någon annan IM-motor än den som installeras automatiskt när du installerar ett språk, kan du <span class="link"><a href="addremove-install.html" title="Installera fler program">installera</a></span> valfri IBus eller Fcitx IM-motor separat.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="keyboard.html" title="Tangentbord">Tangentbord</a><span class="desc"> — <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">Indatakällor</a></span>, <span class="link"><a href="keyboard-cursor-blink.html" title="Gör att tangentbordsmarkören blinkar">blinkande markör</a></span>, <span class="link"><a href="windows-key.html" title='Vad är "Superknappen"?'>supertangent</a></span>, <span class="link"><a href="a11y.html#mobility" title="Rörelsehinder">tangentbordsåtkomst</a></span>...</span>
</li>
<li class="links "><a href="prefs-language.html#textentry" title="Textinmatning">Textinmatning</a></li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="tips-specialchars.html" title="Skriv speciella tecken">Skriv speciella tecken</a><span class="desc"> — Skriv tecken som inte finns på ditt tangentbord, inklusive andra alfabet, matematiska symboler, och dingbats.</span>
</li>
<li class="links ">
<a href="keyboard-shortcuts-set.html" title="Ställ in tangentbordsgenvägar">Ställ in tangentbordsgenvägar</a><span class="desc"> — Definiera eller ändra snabbtangenter i inställningarna för <span class="gui">Tangentbord</span>.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
