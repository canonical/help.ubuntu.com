<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vilka program använder sig av nätkonton?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="accounts.html" title="Nätkonton">Nätkonton</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Vilka program använder sig av nätkonton?</span></h1></div>
<div class="region">
<div class="contents"><p class="p"><span class="app">Nätkonton</span> kan användas av externa program för att automatiskt konfigurera dem.</p></div>
<div id="accounts-google-services" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Med ett Google-konto</span></h2></div>
<div class="region"><div class="contents"><div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p"><span class="app">Evolution</span>, e-postprogrammet. Ditt e-postkonto kommer att läggas till automatiskt i <span class="app">Evolution</span>, så det kan hämta din post, ge dig tillgång till dina kontakter och visa dina kalenderobjekt i din Google-agenda.</p></li>
<li class="list"><p class="p"><span class="app">Empathy</span>, snabbmeddelandeprogrammet. Ditt nätkonto kommer att läggas till och du kommer att kunna kommunicera med dina vänner.</p></li>
<li class="list"><p class="p"><span class="app">Kontakter</span>, kommer att låta dig se och redigera dina kontakter.</p></li>
<li class="list"><p class="p"><span class="app">Dokument</span> kan komma åt dina dokument som lagrats på nätet och visa dem.</p></li>
</ul></div></div></div></div></div>
</div></div>
<div id="accounts-windows-services" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Med Windows Live, Facebook eller Twitter-konton</span></h2></div>
<div class="region"><div class="contents"><p class="p"><span class="app">Empathy</span> kan använda dessa konton för att ansluta till och chatta med dina kontakter, vänner, och följare.</p></div></div>
</div></div>
<div id="account-windows-skydrive" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Med ett SkyDrive-konto</span></h2></div>
<div class="region"><div class="contents"><p class="p"><span class="app">Dokument</span> kan komma åt dina nätdokument i Microsoft SkyDrive och visa dem.</p></div></div>
</div></div>
<div id="account-exchange" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Med ett Exchange-konto</span></h2></div>
<div class="region"><div class="contents"><p class="p">När du har skapat ett Exchange-konto kan <span class="app">Evolution</span> börja hämta e-post från detta konto.</p></div></div>
</div></div>
<div id="accounts-ownCloud" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Med ett ownCloud-konto</span></h2></div>
<div class="region"><div class="contents">
<p class="p">När ett ownCloud-konto är inställt kan <span class="app">Evolution</span> nå och redigera kontakter och kalenderbokningar.</p>
<p class="p"><span class="app">Filer</span> och andra program kommer att kunna lista och nå dina nätfiler sparade i ownCloud-installationen.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="accounts.html" title="Nätkonton">Nätkonton</a><span class="desc"> — <span class="link"><a href="accounts-add.html" title="Lägg till ett konto">Lägg till kontakter, </a></span> <span class="link"><a href="accounts-remove.html" title="Ta bort ett konto">Ta bort konton, </a></span> <span class="link"><a href="accounts-disable-service.html" title="Avaktivera kontotjänster">Avaktivera tjänster</a></span></span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
