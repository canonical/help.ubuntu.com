<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Använda fönster och arbetsytor</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 18.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="getting-started.html.sv" title="Komma igång">Börja med GNOME</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="gs-switch-tasks.html.sv" title="Växla uppgifter">Föregående</a><a class="nextlinks-next" href="gs-use-system-search.html.sv" title="Använd systemsökning">Nästa</a>
</div>
<div class="hgroup"><h1 class="title"><span class="title">Använda fönster och arbetsytor</span></h1></div>
<div class="region">
<div class="contents"><div class="ui-tile ">
<a href="figures/gnome-windows-and-workspaces.webm" class="ui-overlay"><span class="ui-tile-img" style="width: 812px; height: 452px;"><img src="gs-thumb-windows-and-workspaces.svg" width="812" height="452"></span></a><div class="ui-overlay"><div class="inner">
<a href="#" class="ui-overlay-close" title="Stäng">⨯</a><div class="contents"><div class="media media-video"><div class="inner">
<video src="figures/gnome-windows-and-workspaces.webm" preload="auto" controls="controls" class="media media-block" height="394" width="700" data-play-label="Spela upp" data-pause-label="Paus"></video><div class="media-ttml">
<div class="media-ttml-node media-ttml-div" data-ttml-begin="1" data-ttml-end="5"><div class="media-ttml-node media-ttml-p" data-ttml-begin="1" data-ttml-end="5">Fönster och arbetsytor</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="6" data-ttml-end="10"><div class="media-ttml-node media-ttml-p" data-ttml-begin="6" data-ttml-end="10">För att maximera ett fönster, fånga fönstrets namnlist och dra det till toppen på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="10" data-ttml-end="13"><div class="media-ttml-node media-ttml-p" data-ttml-begin="10" data-ttml-end="13">När skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="14" data-ttml-end="20"><div class="media-ttml-node media-ttml-p" data-ttml-begin="14" data-ttml-end="20">För att avmaximera ett fönster, fånga fönstrets namnlist och dra det bort ifrån kanterna på skärmen.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="25" data-ttml-end="29"><div class="media-ttml-node media-ttml-p" data-ttml-begin="25" data-ttml-end="29">Du kan också klicka på namnlisten för att dra bort fönstret och avmaximera det.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="34" data-ttml-end="38"><div class="media-ttml-node media-ttml-p" data-ttml-begin="34" data-ttml-end="38">För att maximera ett fönster längs skärmens vänstra sida, fånga fönstrets namnlist och dra det åt vänster.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="38" data-ttml-end="40"><div class="media-ttml-node media-ttml-p" data-ttml-begin="38" data-ttml-end="40">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="41" data-ttml-end="44"><div class="media-ttml-node media-ttml-p" data-ttml-begin="41" data-ttml-end="44">För att maximera ett fönster längs skärmens högra sida, fånga fönstrets namnlist och dra det åt höger.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="44" data-ttml-end="48"><div class="media-ttml-node media-ttml-p" data-ttml-begin="44" data-ttml-end="48">När halva skärmen är markerad, släpp fönstret.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="54" data-ttml-end="60"><div class="media-ttml-node media-ttml-p" data-ttml-begin="54" data-ttml-end="60">För att maximera ett fönster med tangentbordet, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>↑</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="61" data-ttml-end="66"><div class="media-ttml-node media-ttml-p" data-ttml-begin="61" data-ttml-end="66">För att återställa fönstret till dess avmaximerade storlek, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>↓</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="66" data-ttml-end="73"><div class="media-ttml-node media-ttml-p" data-ttml-begin="66" data-ttml-end="73">För att maximera ett fönster längs den högra sidan på skärmen, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>→</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="76" data-ttml-end="82"><div class="media-ttml-node media-ttml-p" data-ttml-begin="76" data-ttml-end="82">För att maximera ett fönster längs den vänstra sidan på skärmen, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>←</kbd></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="83" data-ttml-end="89"><div class="media-ttml-node media-ttml-p" data-ttml-begin="83" data-ttml-end="89">För att flytta till en arbetsyta som är under den nuvarande arbetsytan, tryck på <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super </kbd></a></span>+<span class="key"><kbd>Page Down</kbd></span></span>.</div></div>
<div class="media-ttml-node media-ttml-div" data-ttml-begin="90" data-ttml-end="97"><div class="media-ttml-node media-ttml-p" data-ttml-begin="90" data-ttml-end="97">För att flytta till en arbetsyta som är ovanför den nuvarande arbetsytan, tryck på <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super </kbd></a></span>+<span class="key"><kbd>Page Up</kbd></span></span>.</div></div>
</div>
</div></div></div>
</div></div>
</div></div>
<div id="use-workspaces-and-windows-maximize" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Maximera och avmaximera fönster</span></h2></div>
<div class="region"><div class="contents">
<p class="p"></p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">För att maximera ett fönster så att det tar upp allt utrymme på ditt skrivbord, fånga fönstrets namnlist och dra det till toppen av skärmen.</p></li>
<li class="steps"><p class="p">När skärmen är markerad, släpp fönstret för att maximera det.</p></li>
<li class="steps"><p class="p">För att återställa ett fönster till dess avmaximerade storlek, fånga fönstrets namnlist och dra det bort från skärmens kanter.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="use-workspaces-and-windows-tile" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Lägg fönster sida-vid-sida</span></h2></div>
<div class="region"><div class="contents">
<p class="p"></p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">För att maximera ett fönster längs en sida av skärmen, fånga fönstrets namnlist och dra det till vänster eller höger sida av skärmen.</p></li>
<li class="steps"><p class="p">När hälften av skärmen är markerad, släpp fönstret för att maximera det längs den valda sidan av skärmen.</p></li>
<li class="steps"><p class="p">För att maximera två fönster sida-vid-sida, fånga namnlisten på det andra fönstret och dra det till den andra sidan av skärmen.</p></li>
<li class="steps"><p class="p">När hälften av skärmen är markerad, släpp fönstret för att maximera det längs den andra sidan av skärmen.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="use-workspaces-and-windows-maximize-keyboard" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Maximera och avmaximera fönster från tangentbordet</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">För att maximera ett fönster med tangentbordet, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>↑</kbd></span>.</p></li>
<li class="steps"><p class="p">För att avmaximera ett fönster genom att använda tangentbordet, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>↓</kbd></span>.</p></li>
</ol></div></div></div></div></div>
</div></div>
<div id="use-workspaces-and-windows-tile-keyboard" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Lägg fönster sida-vid-sida från tangentbordet</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">För att maximera ett fönster längs den högra sidan på skärmen, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>→</kbd></span>.</p></li>
<li class="steps"><p class="p">För att maximera ett fönster längs den vänstra sidan på skärmen, håll ner <span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span> och tryck på <span class="key"><kbd>←</kbd></span>.</p></li>
</ol></div></div></div></div></div>
</div></div>
<div id="use-workspaces-and-windows-workspaces-keyboard" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Växla arbetsytor från tangentbordet</span></h2></div>
<div class="region"><div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">För att flytta till en arbetsyta som är nedanför den aktuella arbetsytan, tryck på <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>+<span class="key"><kbd>Page Down</kbd></span></span>.</p></li>
<li class="steps"><p class="p">För att flytta till en arbetsyta som är ovanför den aktuella arbetsytan, tryck på <span class="keyseq"><span class="key"><a href="help:gnome-help/keyboard-key-super" title="help:gnome-help/keyboard-key-super"><kbd>Super</kbd></a></span>+<span class="key"><kbd>Page Up</kbd></span></span>.</p></li>
</ol></div></div></div></div></div>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="gs-switch-tasks.html.sv" title="Växla uppgifter">Föregående</a><a class="nextlinks-next" href="gs-use-system-search.html.sv" title="Använd systemsökning">Nästa</a>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="getting-started.html.sv" title="Komma igång">Börja med GNOME</a><span class="desc"> — Är GNOME nytt för dig? Lär dig hur du använder det.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="shell-windows-switching.html.sv" title="Växla mellan fönster">Växla mellan fönster</a><span class="desc"> — Tryck <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tabb</kbd></span></span>.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
