<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Why won't DVDs play?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="media.html" title="Ljud, video och bilder">Ljud, video och bilder</a> › <a class="trail" href="media.html#videos" title="Videor och videokameror">Videor</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Why won't DVDs play?</span></h1></div>
<div class="region">
<div class="contents"><p class="p">If you insert a DVD into your computer and it doesn't play, you may not
 have the right DVD <span class="em">codecs</span> installed, or the DVD might be from a
 different <span class="em">region</span>.</p></div>
<div id="codecs" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Installing the right codecs for DVD playback</span></h2></div>
<div class="region"><div class="contents">
<p class="p">In order to play DVDs, you need to have the right <span class="em">codecs</span> installed.
 A codec is a piece of software that allows applications to read a video or
 audio format. If you try to play a DVD and don't have the right codecs installed, the
Movie Player should tell you about this and offer to install them for you.</p>
<p class="p">DVDs are also <span class="em">copy-protected</span> using a system called CSS. This
 prevents you from copying DVDs, but it also prevents you from playing them
 unless you have <span class="link"><a href="video-dvd-restricted.html" title="How do I enable restricted codecs to play DVDs?">extra software</a></span> to handle the copy protection.</p>
</div></div>
</div></div>
<div id="region" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Checking the DVD region</span></h2></div>
<div class="region"><div class="contents">
<p class="p">DVDs have a <span class="em">region code</span>, which tells you in which region of the
 world they are allowed to be played. If the region of your computer's DVD
 player doesn't match the region of the DVD you are trying to play, you won't be
 able to play the DVD. For example, if you have a Region 1 DVD player, you will
 only be allowed to play DVDs from North America.</p>
<p class="p">It is often possible to change the region used by your DVD player, but it
 can only be done a few times before it locks into one region permanently. To
 change the DVD region of your computer's DVD player, use
 <span class="link"><a href="https://apps.ubuntu.com/cat/applications/regionset" title="https://apps.ubuntu.com/cat/applications/regionset">regionset</a></span>.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="media.html#videos" title="Videor och videokameror">Videor</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="video-dvd-restricted.html" title="How do I enable restricted codecs to play DVDs?">How do I enable restricted codecs to play DVDs?</a><span class="desc"> — Most commercial DVDs are encrypted and will not play without decryption software.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
