<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Social networking from the desktop</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-chat.html" title="Chatt &amp; sociala medier">Chatt &amp; sociala medier</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Social networking from the desktop</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">
    With Ubuntu you can post to your favorite social networking sites from your
    desktop. Ubuntu uses the <span class="app">Friends</span> scope to allow you to
    organize your social networking sites in one place, and to post updates
    from the <span class="gui">Me Menu</span> without opening any website.
  </p>
<p class="p"> 
    To set up your social networking accounts:
  </p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">
      Open the <span class="link"><a href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen">System menu</a></span> on the right hand side of the menu bar and select "System Settings...".
    </p></li>
<li class="steps"><p class="p">
      Choose <span class="gui">Online accounts</span>
    </p></li>
<li class="steps"><p class="p">
      Choose the social networking site you want to set up and click <span class="gui">Add Account...</span>
    </p></li>
<li class="steps"><p class="p">
      Click <span class="gui">Authorize</span> and insert your account settings for that site,
      and follow the instructions
    </p></li>
</ol></div></div></div>
<p class="p">
    You can now view your social networking messages from the <span class="link"><a href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen">
    Messaging menu</a></span> 
    on the right hand side of the menu bar, in the <span class="gui">Broadcast</span> section.
    Click on any of the items in that section to open <span class="gui">Friends</span> scope
    and to read or post messages to your social network.
  </p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-chat.html" title="Chatt &amp; sociala medier">Chatt &amp; sociala medier</a><span class="desc"> — 
      <span class="link"><a href="net-chat-empathy.html" title="Snabbmeddelanden på Ubuntu">Chat on any network using <span class="app">Empathy</span></a></span>,
      <span class="link"><a href="net-chat-video.html" title="Video calls">make video calls</a></span>,
      <span class="link"><a href="net-chat-skype.html" title="Hur använder jag Skype på Ubuntu?">install skype</a></span>,
      <span class="link"><a href="net-chat-social.html" title="Social networking from the desktop">social networking apps</a></span>
    </span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
