<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Få ut det mesta ur din bärbara dators batteri</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="power.html" title="På/av &amp; batteri">På/av &amp; batteri</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="power.html" title="På/av &amp; batteri">På/av &amp; batteri</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Få ut det mesta ur din bärbara dators batteri</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Efterhand som batterier åldras blir de sämre på att spara laddning och deras kapacitet minskar gradvis. Det finns ett par tekniker som du kan använda för att förlänga deras användbara livslängd, även om du inte bör förvänta dig en stor skillnad.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list" style="list-style-type:disc">
<li class="list"><p class="p">Låt inte batteriet laddas ur helt. Ladda alltid <span class="em">innan</span> batteriet blir väldigt lågt, även om de flesta batteri har inbyggda skyddsmekanismer för att förhindra att batteriet blir allt för lågt. Att ladda när det bara är delvis urladdat är mer effektivt, men att ladda när det bara är lite urladdat är värre för batteriet.</p></li>
<li class="list"><p class="p">Värme har en skadlig effekt på batteriets laddningseffektivitet. Låt inte batteriet blir varmare än nödvändigt.</p></li>
<li class="list"><p class="p">Batteriet åldras även om du låter dem ligga. Det är bara en liten vinst att köpa ett ersättningsbatteri samtidigt som du köper originalbatteriet - köp alltid ersättningsbatteriet när du behöver dem.</p></li>
</ul></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Detta råd gäller speciellt för Litiumjonbatterier (Li-Ion) vilket är den vanligaste typen. Andra typer av batteriet kan dra fördel av annan behandling.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="power.html" title="På/av &amp; batteri">På/av &amp; batteri</a><span class="desc"> — <span class="link"><a href="power-suspend.html" title="Vad händer när jag försätter min dator i vänteläge?">Vänteläge</a></span>, <span class="link"><a href="power-batterylife.html" title="Använd mindre ström och förbättra batteridriftstiden">spara ström</a></span>, <span class="link"><a href="shell-exit.html#shutdown" title="Stäng av eller starta om">stäng av</a></span>, <span class="link"><a href="power-whydim.html" title="Varför tonas min skärm ner efter ett tag?">mörkare skärm</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="power-batterybroken.html" title="Ett felmeddelande visar att mitt batteri har låg kapacitet">Ett felmeddelande visar att mitt batteri har låg kapacitet</a><span class="desc"> — Ditt batteri är troligtvis inte trasigt; sannolikt är det bara gammalt.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
