<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Hur man skapar en säkerhetskopia</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> › <a class="trail" href="files.html#backup" title="Säkerhetskopiering">Säkerhetskopiering</a> » <a class="trail" href="backup-why.html" title="Säkerhetskopiera dina viktiga filer">Säkerhetskopiering</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Hur man skapar en säkerhetskopia</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Det enklaste sättet att säkerhetskopiera dina filer och inställningar är att låta ett säkerhetskopieringsprogram hantera processen åt dig. Ett antal olika säkerhetskopieringsprogram finns tillgängliga, till exempel <span class="app">Déjà Dup</span>.</p>
<p class="p">Hjälptexten för det kopieringsprogram du väljer kommer vägleda dig genom inställningarna för kopieringen, och hur du återställer dina data.</p>
<p class="p">Ett alternativ är att <span class="link"><a href="files-copy.html" title="Kopiera eller flytta filer och mappar">kopiera dina filer</a></span> till en tillförlitlig plats, exempelvis en extern hårddisk, en annan dator på nätverket eller en USB-enhet. Dina <span class="link"><a href="backup-thinkabout.html" title="Var kan jag hitta filerna jag vill säkerhetskopiera?">personliga filer</a></span> och inställningar finns vanligtvis i din Hemmapp, så du kan kopiera dem därifrån.</p>
<p class="p">Mängden data du kan säkerhetskopiera begränsas av lagringsenhetens utrymme. Om du har tillräckligt mycket utrymme på din säkerhetskopieringsenhet är det bäst att kopiera hela Hemmappen, med följande undantag:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Filer som redan finns säkerhetskopierade någon annanstans, så som på en cd, dvd eller annan flyttbar media.</p></li>
<li class="list"><p class="p">Filer som du kan återställa enkelt. Om du till exempel är en programmerare behöver du inte säkerhetskopiera filer som skapas när du kompilerar dina program. Försäkra dig istället om att du säkerhetskopierar källkodsfilerna.</p></li>
<li class="list"><p class="p">Filer i Papperskorgen. Din Papperskorgsmapp hittar du i <span class="file">~/.local/share/Trash</span>.</p></li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="backup-why.html" title="Säkerhetskopiera dina viktiga filer">Säkerhetskopiera dina viktiga filer</a><span class="desc"> — Varför, vad, var och hur man säkerhetskopierar.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
