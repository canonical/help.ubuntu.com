<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Anslut din dator till en Bluetooth-enhet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="bluetooth.html" title="Bluetooth">Bluetooth</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Anslut din dator till en Bluetooth-enhet</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Innan du kan använda en Bluetooth-enhet som en mus eller ett par hörlurar, måste du först ansluta din dator till enheten. Detta kallas också att <span class="em">para</span> Bluetooth-enheterna.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Bluetooth</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Bluetooth</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Försäkra dig om att Bluetooth är aktiverat: knappen på titelraden ska vara ställd till <span class="gui">PÅ</span>. Med panelen öppen och knappen <span class="gui">PÅ</span>, så kommer din dator att börja söka efter enheter.</p></li>
<li class="steps"><p class="p">Gör din andra Bluetooth-enhet <span class="link"><a href="bluetooth-visibility.html" title="Vad är Bluetooth-synlighet?">detekterbar eller synlig</a></span> och placera den inom 5-10 meter från din dator.</p></li>
<li class="steps"><p class="p">Klicka på enheten i listan <span class="gui">Enheter</span>. Panelen för den enheten kommer att öppnas.</p></li>
<li class="steps">
<p class="p">Om det behövs, bekräfta PIN-koden på din andra enhet. Enheten bör visa PIN-koden du ser på din datorskärm. Bekräfta PIN-koden på enheten (du kan behöva klicka på <span class="gui">Para</span> eller <span class="gui">Bekräfta</span>), klicka sedan på <span class="gui">Bekräfta</span> på datorn.</p>
<p class="p">Du måste avsluta din inmatning inom cirka 20 sekunder för de flesta enheter, annars kommer anslutningen inte att slutföras. Om det händer, gå tillbaka till enhetslistan och börja om igen.</p>
</li>
<li class="steps"><p class="p">Posten för enheten i listan <span class="gui">Enheter</span> kommer att visa statusen <span class="gui">Ansluten</span>.</p></li>
<li class="steps"><p class="p">För att redigera enheten, klicka på den i listan <span class="gui">Enheter</span>. Du kommer att se en panel specifik för den enheten. Den kan visa ytterligare alternativ för den typ av enhet som du ansluter.</p></li>
<li class="steps"><p class="p">Stäng panelen när du har ändrat inställningarna.</p></li>
</ol></div></div></div>
<div class="media media-image floatend"><div class="inner"><img src="figures/bluetooth-menu.png" class="media media-block" alt="Bluetooth-ikonen i systemraden"></div></div>
<p class="p">När en eller flera Bluetooth-enheter är anslutna kommer Bluetooth-ikonen att visas i systemstatusområdet.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="bluetooth.html" title="Bluetooth">Bluetooth</a><span class="desc"> — <span class="link"><a href="bluetooth-connect-device.html" title="Anslut din dator till en Bluetooth-enhet">Anslut</a></span>, <span class="link"><a href="bluetooth-send-file.html" title="Skicka filer till en Bluetooth-enhet">skicka filer</a></span>, <span class="link"><a href="bluetooth-turn-on-off.html" title="Aktivera eller inaktivera Bluetooth">aktivera och inaktivera</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="bluetooth-remove-connection.html" title="Koppla ifrån en Bluetooth-enhet">Koppla ifrån en Bluetooth-enhet</a><span class="desc"> — Ta bort en enhet från listan över Bluetooth-enheter.</span>
</li>
<li class="links ">
<a href="sharing-bluetooth.html" title="Styr delning över Bluetooth">Styr delning över Bluetooth</a><span class="desc"> — Låt filer skickas till din dator över Bluetooth.</span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
