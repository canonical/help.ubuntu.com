<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Bläddra bland filer på en server eller nätverksdelning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="sharing.html" title="Sharing">Sharing</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Bläddra bland filer på en server eller nätverksdelning</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan ansluta till en server eller nätverksdelning för att bläddra bland och visa filer på den servern, precis som om de fanns på din egen dator. Detta är ett bekvämt sätt att ladda ner eller upp filer till internet, eller för att dela filer med andra personer i ditt lokala nätverk.</p>
<p class="p">För att bläddra bland filer i nätverket, öppna programmet <span class="app">Filer</span> från <span class="gui">Dash</span>, och klicka på <span class="gui">Bläddra nätverk</span> i sidoraden. Filhanteraren kommer leta upp datorer i ditt lokala nätverk som signalerar att de kan dela ut sina filer. Om du vill ansluta till en server på internet, eller om du inte ser den dator du letar efter, kan du manuellt ansluta till en server genom att skriva in dess internet-/nätverksadress.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Anslut till en filserver</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">I filhanteraren, klicka på <span class="gui">Filer</span> i menyraden och välj <span class="gui">Anslut till server</span> från programmenyn.</p></li>
<li class="steps">
<p class="p">Skriv serverns adress, i form av en <span class="link"><a href="#urls" title="Skriva URL:er">URL</a></span>. Detaljerad information för URL:er som stöds finns i <span class="link"><a href="#types" title="Typ av servrar">listan nedanför</a></span>.</p>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du har anslutit till servern tidigare kan du klicka på den i listan över <span class="gui">Senaste servrar</span>.</p></div></div></div></div>
</li>
<li class="steps"><p class="p">Klicka på <span class="gui">Anslut</span>. Ett nytt fönster kommer öppnas som visar dig filerna som finns på servern. Du kan bläddra bland filerna precis som om de fanns på din egen dator. Servern kommer också läggas till i sidoraden så att du snabbt kan komma åt den vid ett senare tillfälle</p></li>
</ol></div>
</div></div>
</div>
<div id="urls" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Skriva URL:er</span></h2></div>
<div class="region"><div class="contents">
<p class="p">En <span class="em">URL</span>, eller <span class="em">uniform resource locator</span>, är en typ av adress som hänvisar till en plats eller fil på ett nätverk. Adressen är formaterad så här:</p>
<div class="example"><p class="p"><span class="sys">schema://servernamn.exempel.se/mapp</span></p></div>
<p class="p"><span class="em">Schemat</span> anger vilket protokoll servern använder. <span class="em">Exempel.se</span>-delen av adressen kallas <span class="em">domännamnet</span>. Om ett användarnamn krävs, skrivs det innan servernamnet:</p>
<div class="example"><p class="p"><span class="sys">schema://användarnamn@servernamn.exempel.se/mapp</span></p></div>
<p class="p">Vissa scheman kräver att ett portnummer anges. Skriv det efter domännamnet:</p>
<div class="example"><p class="p"><span class="sys">schema://servernamn.exempel.se:port/mapp</span></p></div>
<p class="p">Nedanför står specifika exempel för de olika servertyper som hanteras.</p>
</div></div>
</div></div>
<div id="types" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Typ av servrar</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan ansluta till olika typer av servrar. En del servrar är allmänna, och låter vem som helst ansluta. Andra servrar kräver att du loggar in med användarnamn och lösenord.</p>
<p class="p">Du har inte alltid tillstånd att utföra vissa åtgärder på filer på en server. På till exempel allmänna FTP-servrar kommer du sannolikt inte kunna radera filer.</p>
<p class="p">URL:en du skriver beror på det protokoll servern använder för att exportera dess delade filer.</p>
<div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">SSH</dt>
<dd class="terms">
<p class="p">Om du har ett <span class="em">secure shell</span>-konto på en server kan du ansluta med den metoden. Många webbhotell delar ut SSH-konton till sina medlemmar så att de kan ladda upp filer på ett säkert sätt. SSH-servrar kräver alltid att du loggar in.</p>
<p class="p">En typisk SSH-URL ser ut så här:</p>
<div class="example"><p class="p"><span class="sys">ssh://användarnamn@servernamn.exempel.se/mapp</span></p></div>
<p class="p">När du använder SSH är all data du skickar (inklusive ditt lösenord) krypterad, så att andra användare på ditt nätverk inte kan se.</p>
</dd>
<dt class="terms">FTP (med inloggning)</dt>
<dd class="terms">
<p class="p">FTP är ett populärt sätt att dela ut filer på internet. Eftersom datan inte krypteras över FTP erbjuder många servrar nu åtkomst via SSH. Vissa servrar, däremot, tillåter eller kräver fortfarande att du använder FTP för upp- eller nedladdning av filer. FTP-sidor med inloggning låter dig ofta radera och ladda upp filer.</p>
<p class="p">En typisk FTP-URL ser ut så här:</p>
<div class="example"><p class="p"><span class="sys">ftp://användarnamn@ftp.exempel.se/sökväg/</span></p></div>
</dd>
<dt class="terms">Offentlig FTP</dt>
<dd class="terms">
<p class="p">Sidor som låter dig ladda ner filer kommer ibland tillåta offentlig eller anonym FTP-anslutning. Dessa servrar kräver inte användarnamn eller lösenord, och kommer i regel inte låta dig radera eller ladda upp filer.</p>
<p class="p">En typisk anonym FTP-URL ser ut så här:</p>
<div class="example"><p class="p"><span class="sys">ftp://ftp.exempel.se/sökväg/</span></p></div>
<p class="p">Vissa anonyma FTP-sidor kräver att du loggar in med ett offentligt användarnamn och lösenord, eller med ett offentligt användarnamn med din e-postadress som lösenord. Använd metoden <span class="gui">FTP (med inloggning)</span>, och använd inloggningsinformationen som efterfrågas av FTP-sidan.</p>
</dd>
<dt class="terms">Windows-utdelning</dt>
<dd class="terms">
<p class="p">Windows-datorer använder ett slutet protokoll för att dela filer i ett lokalt nätverk. Datorer i ett Windows-nätverk grupperas ibland i <span class="em">domäner</span> för bättre organisation och för att ge bättre åtkomstkontroll. Om du har rätt behörighet på fjärrdatorn du är ansluten till kan du ansluta till en Windows-utdelning från filhanteraren.</p>
<p class="p">En typisk URL till en Windows-utdelning ser ut så här:</p>
<div class="example"><p class="p"><span class="sys">smb://servernamn/Utdelning</span></p></div>
</dd>
<dt class="terms">WebDAV och Säker WebDAV</dt>
<dd class="terms">
<p class="p">WebDAV, som bygger på protokollet HTTP, används ibland för att dela filer på ett lokalt nätverk, och för att lagra filer på internet. Om servern du ansluter till har stöd för säkra anslutningar bör du välja det alternativet. Säker WebDAV använder stark SSL-kryptering, så att andra användare inte kan se ditt lösenord.</p>
<p class="p">En typisk WebDAV-URL ser ut så här:</p>
<div class="example"><p class="p"><span class="sys">http://exempel.värdnamn.se/sökväg</span></p></div>
</dd>
</dl></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li>
<li class="links ">
<a href="sharing.html" title="Sharing">Sharing</a><span class="desc"> — 
      <span class="link"><a href="sharing-desktop.html" title="Share your desktop">Desktop sharing</a></span>,
      <span class="link"><a href="files-share.html" title="Dela ut och överför filer">Share files</a></span>…
    </span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-share.html" title="Dela ut och överför filer">Dela ut och överför filer</a><span class="desc"> — För över filer till dina e-postkontakter från filhanteraren.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
