<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Trådlös anslutning</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Trådlös anslutning</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="net-wireless-connect.html" title="Connect to a wireless network"><span class="title">Connect to a wireless network</span><span class="linkdiv-dash"> — </span><span class="desc">Get on the internet - wirelessly.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-vpn-connect.html" title="Connect to a VPN"><span class="title">Connect to a VPN</span><span class="linkdiv-dash"> — </span><span class="desc">VPNs allow you to connect to a local network over the internet. Learn how to set up a VPN connection.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-hidden.html" title="Connect to a hidden wireless network"><span class="title">Connect to a hidden wireless network</span><span class="linkdiv-dash"> — </span><span class="desc">Click the <span class="gui">network menu</span> on the menu bar and select <span class="gui">Connect to Hidden Wireless Network</span>.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-adhoc.html" title="Create a wireless hotspot"><span class="title">Create a wireless hotspot</span><span class="linkdiv-dash"> — </span><span class="desc">Use an ad-hoc network to allow other devices to connect to your
    computer and its network connections.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-find.html" title="I can't see my wireless network in the list"><span class="title">I can't see my wireless network in the list</span><span class="linkdiv-dash"> — </span><span class="desc">The wireless could be turned off or broken, there might be too many wireless networks nearby, or you might be out of range.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-noconnection.html" title="I've entered the correct password, but I still can't connect"><span class="title">I've entered the correct password, but I still can't connect</span><span class="linkdiv-dash"> — </span><span class="desc">Double-check the password, try using the pass key instead of the password, turn the wireless card off and on again…</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="net-manual.html" title="Manually set network settings"><span class="title">Manually set network settings</span><span class="linkdiv-dash"> — </span><span class="desc">If network settings don't get assigned automatically, you may have to enter them yourself.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-edit-connection.html" title="Redigera en trådlös anslutning"><span class="title">Redigera en trådlös anslutning</span><span class="linkdiv-dash"> — </span><span class="desc">Learn what the options on the wireless connection editing screen mean.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-airplane.html" title="Turn off wireless (airplane mode)"><span class="title">Turn off wireless (airplane mode)</span><span class="linkdiv-dash"> — </span><span class="desc">Click the network menu on the menu bar and uncheck Enable Wireless.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?"><span class="title">What do WEP and WPA mean?</span><span class="linkdiv-dash"> — </span><span class="desc">WEP and WPA are ways of encrypting data on wireless networks.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-disconnecting.html" title="Why does my wireless network keep disconnecting?"><span class="title">Why does my wireless network keep disconnecting?</span><span class="linkdiv-dash"> — </span><span class="desc">You might have low signal, or the network might not be letting you connect properly.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter"><span class="title">Wireless network troubleshooter</span><span class="linkdiv-dash"> — </span><span class="desc">Identify and fix problems with wireless connections</span></a></div>
</div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a><span class="desc"> — <span class="link"><a href="net-wireless.html" title="Trådlös anslutning">Trådlöst</a></span>, <span class="link"><a href="net-wired.html" title="Trådbunden anslutning">trådbundet</a></span>, <span class="link"><a href="net-problem.html" title="Nätverksproblem">anslutnings-problem</a></span>, <span class="link"><a href="net-browser.html" title="Webbläsare">webbnavigering</a></span>, <span class="link"><a href="net-email.html" title="E-post &amp; e-postmjukvara">e-postkonton</a></span>, <span class="link"><a href="net-chat.html" title="Chatt &amp; sociala medier">snabbmeddelanden</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="net-general.html" title="Networking terms &amp; tips">Networking terms &amp; tips</a><span class="desc"> — 
      <span class="link"><a href="net-findip.html" title="Hitta din IP-adress">Find your IP address</a></span>,
      <span class="link"><a href="net-wireless-wepwpa.html" title="What do WEP and WPA mean?">WEP &amp; WPA security</a></span>,
      <span class="link"><a href="net-macaddress.html" title="What is a MAC address?">MAC addresses</a></span>,
      <span class="link"><a href="net-proxy.html" title="Define proxy settings">proxies</a></span>…
    </span>
</li>
<li class="links ">
<a href="net-problem.html" title="Nätverksproblem">Nätverksproblem</a><span class="desc"> — 
      <span class="link"><a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Troubleshooting wireless connections</a></span>,
      <span class="link"><a href="net-wireless-find.html" title="I can't see my wireless network in the list">finding your wifi network</a></span>…
        </span>
</li>
</ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
