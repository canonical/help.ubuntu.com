<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="500" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-search1.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2">
      <ns0:stop id="stop3964-5-0-1-9-6-6" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop style="stop-color: rgb(39, 62, 93); stop-opacity: 1;" offset="0.81554461" id="stop6610-2-9-0-2-7"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath56767">
      <ns0:path ns2:nodetypes="ccccc" ns1:connector-curvature="0" id="path56769" d="m 228.45991,29.202459 833.57379,0 0,290.286071 c -330.23641,0 -408.68316,175.76954 -833.57379,175.76954 z" style="color:#000000;fill:#babdb6;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-7">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6281-1-9-2" width="3.8250003" height="6.3750005" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6267-1-9-2" width="2.8977277" height="5.21591" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2">
      <ns0:rect style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" id="rect6261-6-6-2" width="1.8762827" height="4.8734746" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath987-2">
      <ns0:circle r="60" cy="236" cx="63.999996" id="circle989-0" style="display:inline;opacity:1;fill:#3584e4;fill-opacity:1;stroke:none;stroke-width:4.28571415;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath987-2-4">
      <ns0:circle r="60" cy="236" cx="63.999996" id="circle989-0-6" style="display:inline;opacity:1;fill:#3584e4;fill-opacity:1;stroke:none;stroke-width:4.28571415;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath987-2-4-1">
      <ns0:circle r="60" cy="236" cx="63.999996" id="circle989-0-6-1" style="display:inline;opacity:1;fill:#3584e4;fill-opacity:1;stroke:none;stroke-width:4.28571415;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="411.52772" ns1:cy="401.55062" ns1:document-units="px" ns1:current-layer="g17515" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="2560" ns1:window-height="1374" ns1:window-x="0" ns1:window-y="27" ns1:window-maximized="1" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="656" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-540)">
    <ns0:g id="g11020" transform="translate(-35,-107.36217)">
      <ns0:path transform="translate(2,453.36217)" d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" ns2:ry="17" ns2:rx="17" ns2:cy="278" ns2:cx="120" id="path11014" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
      <ns0:text id="text11016" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan11018" ns2:role="line" style="font-size:14px;line-height:1.25">1</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g transform="matrix(0.75098334,0,0,0.75098334,-60.56959,579.06944)" style="display:inline" id="g17515" ns1:export-filename="/home/jimmac/gfx/redhat/redhat-ux/Products/RHEL/RHEL7/video-jingles/tex/overview.png" ns1:export-xdpi="90" ns1:export-ydpi="90" clip-path="url(#clipPath56767)">
      <ns0:g ns1:label="view-grid" id="g7362" transform="matrix(4,0,0,4,172,-591)" style="display:inline">
        <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" id="rect7364" width="16" height="16" x="20" y="276" ns1:label="a"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="279" x="23.0623" height="2" width="2.0000002" id="rect13363" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13365" width="2.0000002" height="2" x="27.0623" y="279" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="279" x="31.0623" height="2" width="2.0000002" id="rect13367" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13369" width="2.0000002" height="2" x="23.0623" y="283.01562" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="283.01562" x="27.0623" height="2" width="2.0000002" id="rect13371" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13373" width="2.0000002" height="2" x="31.0623" y="283.01562" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="287" x="23.0623" height="2" width="2.0000002" id="rect13375" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
        <ns0:rect style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect13377" width="2.0000002" height="2" x="27.0623" y="287" rx="0.38461545" ry="0.37878788"/>
        <ns0:rect ry="0.37878788" rx="0.38461545" y="287" x="31.0623" height="2" width="2.0000002" id="rect13379" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      </ns0:g>
      <ns0:path ns2:nodetypes="ccccccc" ns1:connector-curvature="0" id="rect10989-4" d="m 239.06066,57.414214 800.87864,0 0,51.485276 c 0,0 -4.0279,-10.606597 -11.0989,-10.96015 L 249,99 c -4.59619,-0.353553 -9.93934,5.5 -9.93934,5.5 z" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:g transform="translate(11,0)" id="g10976-7">
        <ns0:rect style="color:#000000;fill:none;stroke:#000000;stroke-width:3;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect10923-0" width="800" height="600" x="229" y="58"/>
        <ns0:path id="path10955-1" style="fill:none;stroke:#000000;stroke-width:2.37319922px;stroke-linecap:round;stroke-linejoin:miter;stroke-opacity:1" d="m 1028.199,108.766 c 0,-5.89806 -4.7813,-10.6794 -10.6794,-10.6794 l -777.99931,0 c -5.89809,0 -10.6794,4.78134 -10.6794,10.6794" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
        <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#000000;fill-opacity:1;stroke:none" x="628.8465" y="86.187378" id="text10972-5"><ns0:tspan ns2:role="line" id="tspan10974-5" x="628.8465" y="86.187378" style="font-size:21.26189423px;line-height:1.25">14:30</ns0:tspan></ns0:text>
        <ns0:path ns2:nodetypes="ccc" ns1:connector-curvature="0" d="m 370.5196,96.0866 -129.99931,0 c -5.89809,0 -10.6794,4.78134 -10.6794,10.6794" style="fill:none;stroke:#000000;stroke-width:5;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" id="path17186"/>
        <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="238.05931" y="86.187378" id="text56758"><ns0:tspan ns2:role="line" id="tspan56760" x="238.05931" y="86.187378" style="font-size:21.26189423px;line-height:1.25">Aktiviteter</ns0:tspan></ns0:text>
        <ns0:g transform="matrix(1.3315875,0,0,1.3315875,6.2833653,3.1816863)" id="g12006">
          <ns0:g id="g5525" transform="translate(689,-168)" ns1:label="audio-volume-medium" style="display:inline">
            <ns0:path ns2:nodetypes="ccccccccc" id="path5533" d="m 20,222 2.484375,0 2.968754,-3 0.546871,0.0156 0,11 -0.475297,8.3e-4 L 22.484375,227 20,227 l 0,-5 z" style="color:#bebebe;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" ns1:connector-curvature="0"/>
            <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" id="rect5535" width="16" height="16" x="20" y="217" ns1:label="audio-volume-high"/>
            <ns0:path clip-path="url(#clipPath6279-7-9-7)" ns2:type="arc" style="fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path3718-5" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
            <ns0:path clip-path="url(#clipPath6265-3-4-4)" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" ns2:ry="3.1875" ns2:rx="3.1875" ns2:cy="223.9375" ns2:cx="24.9375" id="path3726-1" style="fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" ns2:type="arc" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
            <ns0:path clip-path="url(#clipPath6259-8-81-2)" ns2:type="arc" style="opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" id="path3728-0" ns2:cx="24.9375" ns2:cy="223.9375" ns2:rx="3.1875" ns2:ry="3.1875" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" ns2:open="true" ns2:start="5.4977871" ns2:end="7.0685835"/>
          </ns0:g>
          <ns0:g transform="translate(689,-639)" ns1:label="system-shutdown" id="g4692-3" style="display:inline">
            <ns0:rect style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" id="rect10837-3-0" y="688" x="40" ry="0.15129246" rx="0.14408804" height="16" width="16"/>
            <ns0:path ns2:open="true" ns2:end="10.471045" ns2:start="5.239857" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" d="m 51.52343,689.95141 c 3.340544,1.94594 4.471097,6.23148 2.52516,9.57202 -1.945936,3.34054 -6.231476,4.4711 -9.57202,2.52516 -3.340544,-1.94594 -4.471097,-6.23148 -2.52516,-9.57202 0.612757,-1.05191 1.489249,-1.92583 2.542951,-2.53549" ns2:ry="7" ns2:rx="7" ns2:cy="696" ns2:cx="48" id="path3869-2" style="color:#000000;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:type="arc"/>
            <ns0:path ns2:nodetypes="cc" id="path4710" d="m 48,689 0,5" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns1:connector-curvature="0"/>
          </ns0:g>
          <ns0:g id="g12661" transform="translate(666.07286,-166.91767)" ns1:label="network-wired" style="display:inline">
            <ns0:rect ns1:label="audio-volume-high" y="217" x="20" height="16" width="16" id="rect12673" style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible"/>
            <ns0:path id="rect12675" transform="translate(80,257)" d="m -55.25,-40 c -0.952203,0 -1.75,0.7978 -1.75,1.75 l 0,4.5 c 0,0.9522 0.797797,1.75 1.75,1.75 l 0.125,0 -0.78125,1.5625 -0.71875,1.4375 1.625,0 6,0 1.625,0 -0.71875,-1.4375 L -48.875,-32 l 0.125,0 c 0.952203,0 1.75,-0.7978 1.75,-1.75 l 0,-4.5 c 0,-0.9522 -0.797797,-1.75 -1.75,-1.75 l -6.5,0 z m 0.25,2 6,0 0,4 -6,0 0,-4 z" style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#bebebe;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans" ns1:connector-curvature="0"/>
            <ns0:path style="color:#bebebe;fill:none;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible" d="m 88,196 0,4" id="path12679" transform="translate(-60.0003,30)" ns1:connector-curvature="0"/>
            <ns0:path style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:2;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible" d="m 21.99975,231 12,0" id="path12681" ns1:connector-curvature="0"/>
          </ns0:g>
          <ns0:path ns2:nodetypes="cccc" ns1:connector-curvature="0" id="rect12003" d="m 759.10724,57.4163 -3.74999,3.750004 -3.75001,-3.750005 z" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate"/>
        </ns0:g>
      </ns0:g>
      <ns0:rect ry="24.20339" rx="24.20339" y="121.79661" x="488.77966" height="48.40678" width="290.44067" id="rect11062-3" style="color:#000000;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:3;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:path transform="matrix(2.6034636,0,0,2.6005055,-53.490592,-862.05263)" d="m 311,386.5 c 0,1.933 -1.567,3.5 -3.5,3.5 -1.933,0 -3.5,-1.567 -3.5,-3.5 0,-1.933 1.567,-3.5 3.5,-3.5 1.933,0 3.5,1.567 3.5,3.5 z" ns2:ry="3.5" ns2:rx="3.5" ns2:cy="386.5" ns2:cx="307.5" id="path27918" style="color:#000000;fill:none;stroke:#000000;stroke-width:1.55467153;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns2:type="arc"/>
      <ns0:path ns2:nodetypes="cc" id="path27941" d="m 754.16168,150.12192 8.09967,8.09046" style="color:#000000;fill:none;stroke:#000000;stroke-width:4.04523087;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" ns1:connector-curvature="0"/>
      <ns0:rect style="opacity:0.70638272;color:#000000;fill:none;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" id="rect1431" width="32.361851" height="32.361847" x="733.91248" y="129.89575"/>
      <ns0:path ns2:nodetypes="cssssc" ns1:connector-curvature="0" id="rect17188" d="m 239.70338,191.5 75.59324,0 c 6.76067,0 12.20338,5.44271 12.20338,12.20338 l 0,371.59324 c 0,6.76067 -5.44271,12.20338 -12.20338,12.20338 l -75.59324,0" style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-linecap:square;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new"/>
      <ns0:g style="display:inline" id="g6180" transform="matrix(0.48410848,0,0,0.48410848,484.01337,-3.4388029)">
        <ns0:g style="display:inline;stroke-width:0.93333334;enable-background:new" transform="matrix(0.26785714,0,0,0.26785714,-482.48304,489.73394)" id="g912-6">
          <ns0:circle r="224" cy="43.999989" cx="256" id="circle1036" style="display:inline;opacity:1;fill:#000000;fill-opacity:1;stroke:#000000;stroke-width:14.9333334;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
        </ns0:g>
        <ns0:path ns2:nodetypes="ccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccccc" ns1:connector-curvature="0" id="path991" d="m 38,176 v 4 l 10,8 v 8 l 8,8 h 4 v -4 l 6,-6 v -4 l 4,-4 v -10 z m -4,16 H 4 c 0,0 0.5090211,40.4419 0,40 l 20,18 v -6 l -4,-4 6,-6 h 4 l 4,4 0.12494,-8.4018 L 40,224 h 4 v -4 l 4,-4 v -6 L 43.727619,206.12499 34,206 v 8 h -4 l -4,-4 v -4 l 6,-6 h 6 v -4 z m 60,2 -6,6 v 4 h 6 v -2.14287 h 4 v 4.26786 L 96,208 H 86 v 4 h -4 v 6 h -8 v 8 h 10 v -4 h 8 v 2 l 4,4 h 2 v -2 l -2,-2 v -2 h 4 l 6,6 h 6 v 2 l -2,2 h -4 l 18,18 V 194 H 96 Z m 12,38 H 94 l -2,-2 H 78 l -8,8 v 8 l 8,8 h 6 l 4,4 v 2 l 2,2 v 12 l 14,14 h 8 v -30 l 4,-4 v -8 l -10,-10 z m -2,-12 h 4 l 6,6 h -4 z m -74,28 -4,4 v 10 l 8.12494,8.14285 L 34,296 h 8 v -8 l 6,-6 v -4 l 6,-6 v -4 l 4,-4 v -8 l -4,-4 h -8 l -4,-4 z" clip-path="url(#clipPath987-2-4-1)" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.01129821px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:accumulate" transform="matrix(0.96464464,0,0,0.96464464,-475.64889,273.86349)"/>
        <ns0:g transform="matrix(0.33027944,0,0,0.33027944,-722.51179,363.54416)" id="g6008" style="display:inline;opacity:1;stroke:#000000;enable-background:new">
          <ns0:circle r="36.270779" cy="372.21783" cx="883.60425" id="path3066-4" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:16.92636299;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
          <ns0:circle r="68.971695" cy="372.2179" cx="883.60431" id="path3941-2" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:11.69271851;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
          <ns0:circle r="103.1213" cy="372.21796" cx="883.60437" id="path3943-0" style="color:#000000;display:inline;overflow:visible;visibility:visible;opacity:0.66763006;fill:none;stroke:#000000;stroke-width:5.99500418;stroke-linecap:butt;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none"/>
        </ns0:g>
        <ns0:g transform="translate(-477.91161,277.51965)" id="g6092" style="display:inline;enable-background:new">
          <ns0:g id="g6087">
            <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#ffffff;fill-opacity:1;fill-rule:evenodd;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:new" ns2:nodetypes="cccssccc" id="path3970-7-4" d="m 47.589745,209.314 -47.7665216,46.36163 21.7759096,0.70244 c 0,0 -9.131831,18.96611 -9.131831,18.96611 -2.8097966,8.42939 9.834282,11.59041 11.941628,5.26838 0,0 8.42939,-18.96612 8.42939,-18.96612 l 15.453872,16.50755 z" ns1:connector-curvature="0"/>
          </ns0:g>
        </ns0:g>
      </ns0:g>
      <ns0:path style="color:#000000;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:sans-serif;font-variant-ligatures:normal;font-variant-position:normal;font-variant-caps:normal;font-variant-numeric:normal;font-variant-alternates:normal;font-feature-settings:normal;text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;text-decoration-style:solid;text-decoration-color:#000000;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-orientation:mixed;dominant-baseline:auto;baseline-shift:baseline;text-anchor:start;white-space:normal;shape-padding:0;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:3.87286782;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:new" d="m 261.56425,290.96321 a 5.8093017,5.8093017 0 0 0 -5.80934,5.80929 5.8093017,5.8093017 0 0 0 3.87289,5.46987 v 31.66186 a 5.8093017,5.8093017 0 0 0 -3.87289,5.46984 5.8093017,5.8093017 0 0 0 5.80934,5.80935 5.8093017,5.8093017 0 0 0 5.02545,-2.90469 h 32.55345 a 5.8093017,5.8093017 0 0 0 5.02259,2.90469 5.8093017,5.8093017 0 0 0 5.80935,-5.80935 5.8093017,5.8093017 0 0 0 -3.87291,-5.46984 v -31.66186 a 5.8093017,5.8093017 0 0 0 3.87291,-5.46987 5.8093017,5.8093017 0 0 0 -5.80935,-5.80929 5.8093017,5.8093017 0 0 0 -5.72136,4.84109 h -31.1531 a 5.8093017,5.8093017 0 0 0 -5.72703,-4.84109 z m 5.02545,8.71396 h 32.55345 a 5.8093017,5.8093017 0 0 0 0.1269,0.22134 l -5.01979,5.0198 a 3.8728679,3.8728679 0 0 0 -1.70288,-0.40009 3.8728679,3.8728679 0 0 0 -3.74431,2.90461 h -11.87291 a 3.8728679,3.8728679 0 0 0 -3.74712,-2.90461 3.8728679,3.8728679 0 0 0 -1.70477,0.39802 l -5.02169,-5.02171 a 5.8093017,5.8093017 0 0 0 0.13343,-0.21772 z m -3.08903,2.73824 5.81683,5.81688 a 3.8728679,3.8728679 0 0 0 -0.005,0.15898 3.8728679,3.8728679 0 0 0 1.93642,3.34996 v 12.66628 a 3.8728679,3.8728679 0 0 0 -1.93642,3.34811 3.8728679,3.8728679 0 0 0 0.39801,1.70478 l -5.02171,5.02168 a 5.8093017,5.8093017 0 0 0 -1.1857,-0.57772 z m 38.72866,0 v 31.48882 a 5.8093017,5.8093017 0 0 0 -1.18946,0.57391 l -5.01978,-5.01982 a 3.8728679,3.8728679 0 0 0 0.40009,-1.70283 3.8728679,3.8728679 0 0 0 -1.93641,-3.35005 v -12.6662 a 3.8728679,3.8728679 0 0 0 1.93641,-3.34811 3.8728679,3.8728679 0 0 0 -0.005,-0.16053 z m -26.49168,8.88039 h 14.25284 a 3.8728679,3.8728679 0 0 0 0.62025,0.4453 v 12.66627 a 3.8728679,3.8728679 0 0 0 -1.80787,2.37986 h -11.87294 a 3.8728679,3.8728679 0 0 0 -1.81068,-2.38179 v -12.6662 a 3.8728679,3.8728679 0 0 0 0.6184,-0.44322 z m 0,19.3643 h 14.25284 a 3.8728679,3.8728679 0 0 0 2.55669,0.96823 3.8728679,3.8728679 0 0 0 0.16053,-0.005 l 5.94168,5.94169 a 5.8093017,5.8093017 0 0 0 -0.20523,0.84154 h -31.1531 a 5.8093017,5.8093017 0 0 0 -0.21357,-0.8387 l 5.94643,-5.94639 a 3.8728679,3.8728679 0 0 0 0.15898,0.005 3.8728679,3.8728679 0 0 0 2.55481,-0.96827 z" id="path1558" ns1:connector-curvature="0"/>
      <ns0:g transform="matrix(0.48410848,0,0,0.48410848,251.70413,280.43344)" style="display:inline;enable-background:new" id="g1207">
        <ns0:rect ry="8.555583" rx="8.555583" y="176.2498" x="16.944288" height="115.50041" width="94.111382" id="rect15435-6" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:4;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
        <ns0:path style="display:inline;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.0119126px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" d="m 525,430.125 c -2.216,0 -4,1.784 -4,4 V 463 h 80 v -28.875 c 0,-2.216 -1.784,-4 -4,-4 z M 521,465 v 30 h 80 v -30 z m 0,32 v 29 c 0,2.216 1.784,4 4,4 h 72 c 2.216,0 4,-1.784 4,-4 v -29 z" transform="translate(-497,-247)" id="rect15441-8" ns1:connector-curvature="0" ns2:nodetypes="ssccsssccccccsssscc"/>
        <ns0:g id="g1088">
          <ns0:path style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.01184966px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" d="m 552,443 c -1.662,0 -3,1.338 -3,3 v 4 1 h 4 0.0312 l -0.0156,-2 H 569 v 2 H 569.0312 573 v -1 -4 c 0,-2 -1.338,-3 -3,-3 z" transform="translate(-497,-247)" id="path26035" ns1:connector-curvature="0"/>
        </ns0:g>
        <ns0:use height="100%" width="100%" transform="translate(0,32)" id="use1090" ns4:href="#g1088" y="0" x="0"/>
        <ns0:use x="0" y="0" ns4:href="#g1088" id="use1092" transform="translate(0,64)" width="100%" height="100%"/>
      </ns0:g>
      <ns0:g style="display:inline" transform="matrix(0.48410848,0,0,0.48410848,-125.4164,778.81367)" id="g16105">
        <ns0:path ns1:connector-curvature="0" id="rect854" d="m 798.33622,-694.6285 c -4.70031,0 -8.48432,3.78401 -8.48432,8.48432 v 10.60536 74.23787 8.48433 c 0,4.70031 3.78401,8.48432 8.48432,8.48432 h 93.32756 c 4.70031,0 8.48432,-3.78401 8.48432,-8.48432 v -8.48433 -74.23787 -10.60536 c 0,-4.70031 -3.78401,-8.48432 -8.48432,-8.48432 z" style="display:inline;opacity:1;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:4;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new"/>
        <ns0:rect style="display:inline;opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.01121096px;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;enable-background:new" id="rect858" width="96" height="87.999969" x="797" y="599.48041" rx="4" ry="3.9999695" transform="scale(1,-1)"/>
        <ns0:g style="display:inline;fill:#ffffff;enable-background:new" transform="translate(779,-877.48042)" id="g866">
          <ns0:path ns1:connector-curvature="0" id="path862" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:medium;line-height:1.25;font-family:'Source Code Pro';-inkscape-font-specification:'Source Code Pro, Bold';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.24999999" d="M 44.012301,210.88755 30,203.27182 V 208 l 9.710724,4.62951 v 0.1422 L 30,218 v 4.72818 l 14.012301,-8.21451 z" ns2:nodetypes="ccccccccc"/>
          <ns0:path ns2:nodetypes="ccccc" ns1:connector-curvature="0" id="path864" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;font-size:medium;line-height:1.25;font-family:'Source Code Pro';-inkscape-font-specification:'Source Code Pro, Bold';font-variant-ligatures:normal;font-variant-caps:normal;font-variant-numeric:normal;font-feature-settings:normal;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:0.24999999" d="m 47.999998,226 2e-6,4 h 16.00001 l -2e-6,-4 z"/>
        </ns0:g>
      </ns0:g>
    </ns0:g>
    <ns0:path style="color:#000000;fill:none;stroke:#000000;stroke-width:1;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:2, 4;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" d="M 720.5,819 C 472.49798,819 438.08578,951 119,951" id="rect56762" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
    <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;fill:#000000;fill-opacity:1;stroke:none" x="323.60797" y="692.51361" id="text57298"><ns0:tspan ns2:role="line" id="tspan57300" x="323.60797" y="692.51361" style="font-size:14px;line-height:1.25">bara skriv</ns0:tspan></ns0:text>
  </ns0:g>
</ns0:svg>
