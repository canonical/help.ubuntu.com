<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ström och batteri</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Ström och batteri</span></h1></div>
<div class="region">
<div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-status.html.sv" title="Kontrollera batteristatus"><span class="title">Kontrollera batteristatus</span><span class="linkdiv-dash"> — </span><span class="desc">Visa status för batteriet och anslutna enheter.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-batterylife.html.sv" title="Använd mindre ström och förbättra batteridriftstiden"><span class="title">Använd mindre ström och förbättra batteridriftstiden</span><span class="linkdiv-dash"> — </span><span class="desc">Tips på hur du reducerar din dators strömförbrukning.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-batteryoptimal.html.sv" title="Få ut det mesta ur din bärbara dators batteri"><span class="title">Få ut det mesta ur din bärbara dators batteri</span><span class="linkdiv-dash"> — </span><span class="desc">Tips så som ”Låt inte batteriet bli för lågt”.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-exit.html.sv" title="Logga ut, stäng av eller växla användare"><span class="title">Logga ut, stäng av eller växla användare</span><span class="linkdiv-dash"> — </span><span class="desc">Lär dig hur du lämnar ditt användarkonto genom att logga ut, växla användare, och så vidare.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-wireless.html.sv" title="Slå av trådlösa teknologier som inte används"><span class="title">Slå av trådlösa teknologier som inte används</span><span class="linkdiv-dash"> — </span><span class="desc">Bluetooth, wi-fi och mobilt bredband kan slås av för att minska batterianvändning.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-suspend.html.sv" title="Vad händer när jag försätter min dator i vänteläge?"><span class="title">Vad händer när jag försätter min dator i vänteläge?</span><span class="linkdiv-dash"> — </span><span class="desc">Vänteläge försätter din dator i ett strömsparläge där den drar mindre ström.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-closelid.html.sv" title="Varför stängs min dator av när jag stänger locket?"><span class="title">Varför stängs min dator av när jag stänger locket?</span><span class="linkdiv-dash"> — </span><span class="desc">Bärbara datorer försätts i strömsparläge när du stänger locket för att spara ström.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-percentage.html.sv" title="Visa batteristatus som en procentsats"><span class="title">Visa batteristatus som en procentsats</span><span class="linkdiv-dash"> — </span><span class="desc">Visa batteriprocent i systemraden.</span></a></div>
</div>
</div></div></div></div></div>
<section id="saving"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Strömsparinställningar</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-autobrightness.html.sv" title="Aktivera automatisk ljusstyrka"><span class="title">Aktivera automatisk ljusstyrka</span><span class="linkdiv-dash"> — </span><span class="desc">Styr automatiskt skärmljusstyrka för att minska batterianvändning.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-autosuspend.html.sv" title="Konfigurera automatiskt vänteläge"><span class="title">Konfigurera automatiskt vänteläge</span><span class="linkdiv-dash"> — </span><span class="desc">Konfigurera din dator att automatiskt gå i vänteläge.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="display-blank.html.sv" title="Ställ in tiden för skärmtömning"><span class="title">Ställ in tiden för skärmtömning</span><span class="linkdiv-dash"> — </span><span class="desc">Ändra tiden till skärmtömning för att spara ström.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-whydim.html.sv" title="Varför tonas min skärm ner efter ett tag?"><span class="title">Varför tonas min skärm ner efter ett tag?</span><span class="linkdiv-dash"> — </span><span class="desc">Skärmen tonas ner när datorn är oanvänd för att spara ström.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-profile.html.sv" title="Välj en strömprofil"><span class="title">Välj en strömprofil</span><span class="linkdiv-dash"> — </span><span class="desc">Balansera prestanda och batterianvändning.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="faq"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Frågor</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-batteryestimate.html.sv" title="Den uppskattade batteridriftstiden är fel"><span class="title">Den uppskattade batteridriftstiden är fel</span><span class="linkdiv-dash"> — </span><span class="desc">Batteridriftstiden som visas när du klickar på <span class="gui">batteriikonen</span> är en uppskattning.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-batterywindows.html.sv" title="Varför har jag mindre batteridriftstid än jag hade i Windows/Mac OS?"><span class="title">Varför har jag mindre batteridriftstid än jag hade i Windows/Mac OS?</span><span class="linkdiv-dash"> — </span><span class="desc">Justeringar från tillverkaren och olika batteridriftsuppskattningar kan vara orsaken till detta problem.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-lowpower.html.sv" title="Varför stängdes min dator av när batteriet gick ner till 10%?"><span class="title">Varför stängdes min dator av när batteriet gick ner till 10%?</span><span class="linkdiv-dash"> — </span><span class="desc">Att låta batteriet laddas ur helt är dåligt för batteriet.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-batteryslow.html.sv" title="Varför är min bärbara dator så långsam när den kör på batteri?"><span class="title">Varför är min bärbara dator så långsam när den kör på batteri?</span><span class="linkdiv-dash"> — </span><span class="desc">Vissa bärbara datorer kör avsiktligt saktare när de kör på batteri.</span></a></div>
</div>
</div></div></div></div></div></div>
</div></section><section id="problems"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Problem</span></h2></div>
<div class="region">
<div class="contents pagewide"><div class="links topiclinks"><div class="inner"><div class="region"><div class="links-twocolumn">
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-constantfan.html.sv" title="Den bärbara datorns fläkt kör alltid"><span class="title">Den bärbara datorns fläkt kör alltid</span><span class="linkdiv-dash"> — </span><span class="desc">Någon kontrollprogramvara för fläkten kan saknas, eller så är din dator varm.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-nowireless.html.sv" title="Jag har inget trådlöst nätverk när jag väcker datorn"><span class="title">Jag har inget trådlöst nätverk när jag väcker datorn</span><span class="linkdiv-dash"> — </span><span class="desc">Vissa trådlösa enheter har problem med att hantera när datorn är i vänteläge och återstartar inte korrekt.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-othercountry.html.sv" title="Kommer min dator att fungera med ett strömaggregat i ett annat land?"><span class="title">Kommer min dator att fungera med ett strömaggregat i ett annat land?</span><span class="linkdiv-dash"> — </span><span class="desc">Din dator kommer att fungera, men du kan komma att behöva en annan strömsladd eller en reseadapter.</span></a></div>
</div>
<div class="links-divs">
<div class="linkdiv "><a class="linkdiv" href="power-hotcomputer.html.sv" title="Min dator blir väldigt varm"><span class="title">Min dator blir väldigt varm</span><span class="linkdiv-dash"> — </span><span class="desc">Datorer blir vanligtvis varma, men om de blir allt för varma kan de överhettas vilket kan skada datorn.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-willnotturnon.html.sv" title="Min dator vill inte starta"><span class="title">Min dator vill inte starta</span><span class="linkdiv-dash"> — </span><span class="desc">Lösa kablar och hårdvaruproblem är möjliga orsaker.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-suspendfail.html.sv" title="Varför återstartar inte min dator efter att jag har försatt den i vänteläge?"><span class="title">Varför återstartar inte min dator efter att jag har försatt den i vänteläge?</span><span class="linkdiv-dash"> — </span><span class="desc">Viss datorhårdvara orsakar problem med vänteläge.</span></a></div>
</div>
</div></div></div></div></div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h3><span class="title">Mer information</span></h3></div>
<div class="region"><ul><li class="links "><a href="hardware.html.sv#problems" title="Vanliga problem">Hårdvaruproblem</a></li></ul></div>
</div></div></div>
</div></section>
</div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — Få GNOME att arbeta för dig, från hårdvarukontroll till sekretessinställningar.</span>
</li>
<li class="links ">
<a href="hardware.html.sv" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a><span class="desc"> — Konfigurera hårdvara och diagnostisera problem, inklusive skrivare, skärmar, diskar med mera.</span>
</li>
</ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
