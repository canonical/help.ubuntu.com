<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Anslut till mobilt bredband</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Anslut till mobilt bredband</span></h1></div>
<div class="region">
<div class="contents">
<p class="p"><span class="em">Mobilt bredband</span> avser en godtycklig typ av internetanslutning som tillhandahålls av en extern enhet, som en 3G USB-sticka eller mobiltelefon med inbyggd HSPA/UMTS/GPRS-dataanslutning. Vissa bärbara datorer har nyligen tillverkats med inbyggda enheter för mobilt bredband.</p>
<p class="p">De flesta enheter för mobilt bredband bör kännas igen automatiskt när du ansluter dem till din dator. Ubuntu kommer be dig ställa in enheten.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Guiden <span class="gui">Ny mobilt bredbandsanslutning</span> kommer öppnas automatiskt när du ansluter enheten.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Framåt</span> och fyll i fälten, inklusive landet där din enhet för mobilt bredband skickades från, nätverksleverantör, och anslutningstyp (exempelvis <span class="em">Kontrakt</span> eller <span class="em">förbetalning</span>).</p></li>
<li class="steps"><p class="p">Ge din anslutning ett namn och klicka på <span class="gui">Verkställ</span>.</p></li>
<li class="steps"><p class="p">Din anslutning kan nu användas. För att ansluta, klicka på <span class="gui">nätverksmenyn</span> i <span class="gui">menyraden</span> och välj din nya anslutning.</p></li>
<li class="steps"><p class="p">För att koppla från, klicka på <span class="gui">nätverksmenyn</span> i menyraden och klicka på <span class="gui">Koppla från</span>.</p></li>
</ol></div></div></div>
<p class="p">Om du inte blir ombedd att ställa in enheten när du ansluter den kan den ändå kännas igen av Ubuntu. I sådana fall kan du lägga till anslutningen manuellt.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Klicka på <span class="link"><a href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen">nätverksmenyn</a></span> i menyraden och välj <span class="gui">Redigera anslutningar...</span></p></li>
<li class="steps"><p class="p">Byt till fliken <span class="gui">Mobilt bredband</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Lägg till</span>.</p></li>
<li class="steps"><p class="p">Detta bör öppna guiden <span class="gui">Ny anslutning via mobilt breband</span>. Fyll i fälten som förut.</p></li>
</ol></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a><span class="desc"> — <span class="link"><a href="net-wireless.html" title="Trådlös anslutning">Trådlöst</a></span>, <span class="link"><a href="net-wired.html" title="Trådbunden anslutning">trådbundet</a></span>, <span class="link"><a href="net-problem.html" title="Nätverksproblem">anslutnings-problem</a></span>, <span class="link"><a href="net-browser.html" title="Webbläsare">webbnavigering</a></span>, <span class="link"><a href="net-email.html" title="E-post &amp; e-postmjukvara">e-postkonton</a></span>, <span class="link"><a href="net-chat.html" title="Chatt &amp; sociala medier">snabbmeddelanden</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
