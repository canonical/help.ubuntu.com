<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Lägg till föräldrakontroller</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 23.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="user-accounts.html.sv" title="Användarkonton">Användare</a> › <a class="trail" href="user-accounts.html.sv#manage" title="Hantera användarkonton">Konton</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Lägg till föräldrakontroller</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Föräldrar kan använda programmet <span class="gui">Föräldrakontroller</span> för att förhindra barn från att komma åt skadligt innehåll.</p>
<p class="p">En systemadministratör kan använda detta program för att:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Begränsa en användares åtkomst till webbläsare och program.</p></li>
<li class="list"><p class="p">Förhindra en användare från att installera program.</p></li>
<li class="list"><p class="p">Endast ge en användare åtkomst till program lämpliga för åldern.</p></li>
</ul></div></div></div>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p"><span class="gui">Föräldrakontroller</span> kräver att program installeras via Flatpak eller Flathub.</p></div></div></div>
</div>
</div>
<section id="restrictwebbrowsers"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Begränsa webbläsare</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p"><span class="gui">Föräldrakontroller</span> låter en administratör inaktivera webbläsaråtkomst för en användare.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Användare</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Användare</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Välj under <span class="gui">Andra användare</span> användaren som du vill tillämpa kontrollerna på.</p></li>
<li class="steps">
<p class="p">Välj fliken <span class="gui">Föräldrakontroller</span>.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Fliken visas endast om <span class="gui">Föräldrakontroller</span> är installerat och aktiverat.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Tryck på <span class="gui">Lås upp</span> i dialogrutan <span class="gui">Behörighet krävs</span>.</p></li>
<li class="steps"><p class="p">Ange ditt lösenord och autentisera för att låsa upp dialogrutan <span class="gui">Föräldrakontroller</span>.</p></li>
<li class="steps"><p class="p">Slå på <span class="gui">Begränsa webbläsare</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></section><section id="restrictapplications"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Begränsa program</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p"><span class="gui">Föräldrakontroller</span> tillhandahåller en lista över program som en administratör kan inaktivera.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Befintliga program (som inte installerats via Flatpak) kommer inte visas i denna lista.</p></div></div></div>
</div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Användare</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Användare</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Välj under <span class="gui">Andra användare</span> användaren som du vill tillämpa kontrollerna på.</p></li>
<li class="steps">
<p class="p">Välj fliken <span class="gui">Föräldrakontroller</span>.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Fliken visas endast om <span class="gui">Föräldrakontroller</span> är installerat och aktiverat.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Tryck på <span class="gui">Lås upp</span> i dialogrutan <span class="gui">Behörighet krävs</span>.</p></li>
<li class="steps"><p class="p">Ange ditt lösenord och autentisera för att låsa upp dialogrutan <span class="gui">Föräldrakontroller</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Begränsa program</span>.</p></li>
<li class="steps"><p class="p">Växla brytaren intill det eller de program du vill begränsa.</p></li>
</ol></div></div></div>
</div></div>
</div></section><section id="restrictapplicationinstallation"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Begränsa installation av program</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p"><span class="gui">Föräldrakontroller</span> låter en administratör neka installationsprivilegier för en användare.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Användare</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Användare</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Välj under <span class="gui">Andra användare</span> användaren som du vill tillämpa kontrollerna på.</p></li>
<li class="steps">
<p class="p">Välj fliken <span class="gui">Föräldrakontroller</span>.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Fliken visas endast om <span class="gui">Föräldrakontroller</span> är installerat och aktiverat.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Tryck på <span class="gui">Lås upp</span> i dialogrutan <span class="gui">Behörighet krävs</span>.</p></li>
<li class="steps"><p class="p">Ange ditt lösenord och autentisera för att låsa upp dialogrutan <span class="gui">Föräldrakontroller</span>.</p></li>
<li class="steps"><p class="p">Slå på brytaren <span class="gui">Begränsa installation av program</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></section><section id="applicationsuitability"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Begränsa program efter åldersgrupp</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Begränsa vilka program som är synliga baserat på deras lämplighet för en viss åldersgrupp.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Användare</span>.</p></li>
<li class="steps"><p class="p">Välj <span class="gui">Användare</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Välj under <span class="gui">Andra användare</span> användaren som du vill tillämpa kontrollerna på.</p></li>
<li class="steps">
<p class="p">Välj fliken <span class="gui">Föräldrakontroller</span>.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Fliken visas endast om <span class="gui">Föräldrakontroller</span> är installerat och aktiverat.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Tryck på <span class="gui">Lås upp</span> i dialogrutan <span class="gui">Behörighet krävs</span>.</p></li>
<li class="steps"><p class="p">Ange ditt lösenord och autentisera för att låsa upp dialogrutan <span class="gui">Föräldrakontroller</span>.</p></li>
<li class="steps"><p class="p">Välj åldersgruppen från rullgardinslistan i <span class="gui">Programmet lämpligt för</span>.</p></li>
</ol></div></div></div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="user-accounts.html.sv#manage" title="Hantera användarkonton">Hantera användarkonton</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
