<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Connect to mobile broadband</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Connect to mobile broadband</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">
      <span class="em">Mobile Broadband</span> refers to any kind of high speed 
      Internet connection which is provided by an external device such as a 
      3G USB stick or mobile phone with built-in HSPA/UMTS/GPRS data 
      connection. Some laptops have recently been produced with mobile 
      broadband devices already inside them.
    </p>
<p class="p">
      Most mobile broadband devices should be recognized automatically when you 
      connect them to your computer. Ubuntu will prompt you to configure the 
      device.
    </p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">
          The <span class="gui">New Mobile Broadband Connection</span> wizard will 
          open automatically when you connect the device.
          </p></li>
<li class="steps"><p class="p">
          Click <span class="gui">Forward</span> and enter your details, 
          including the country where your Mobile Broadband device was issued, 
          the network provider and type of connection (for example, 
          <span class="em">Contract</span> or <span class="em">pre-pay</span>).
          </p></li>
<li class="steps"><p class="p">
          Give your connection a name and click <span class="gui">Apply</span>.
          </p></li>
<li class="steps"><p class="p">
          Your connection is now ready to use. To connect, click the <span class="gui">network 
          menu</span> in the <span class="gui">menu bar</span> and select your new connection.
          </p></li>
<li class="steps"><p class="p">
          To disconnect, click the <span class="gui">network menu</span> in the menu bar and click
          <span class="gui">Disconnect</span>.
          </p></li>
</ol></div></div></div>
<p class="p">
    If you are not prompted to configure the device when you connect it, it 
    may still be recognized by Ubuntu. In such cases you can add the connection 
    manually.
    </p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">
    	  Click the <span class="link"><a href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen">network menu</a></span> in the menu bar 
    	  and select <span class="gui">Edit Connections...</span>
    	  </p></li>
<li class="steps"><p class="p">
    	  Switch to the <span class="gui">Mobile Broadband</span> tab.
    	  </p></li>
<li class="steps"><p class="p">
    	  Click <span class="gui">Add</span>.
    	  </p></li>
<li class="steps"><p class="p">
    	  This should open the <span class="gui">New Mobile Broadband 
    	  Connection</span> wizard. Enter your details as described above.
    	  </p></li>
</ol></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a><span class="desc"> — <span class="link"><a href="net-wireless.html" title="Trådlös anslutning">Trådlöst</a></span>, <span class="link"><a href="net-wired.html" title="Trådbunden anslutning">trådbundet</a></span>, <span class="link"><a href="net-problem.html" title="Nätverksproblem">anslutnings-problem</a></span>, <span class="link"><a href="net-browser.html" title="Webbläsare">webbnavigering</a></span>, <span class="link"><a href="net-email.html" title="E-post &amp; e-postmjukvara">e-postkonton</a></span>, <span class="link"><a href="net-chat.html" title="Chatt &amp; sociala medier">snabbmeddelanden</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
