<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Sök efter filer</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Sök efter filer</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan söka efter filer baserat på namn eller filtyp direkt från filhanteraren. Du kan också spara vanliga sökningar, och de kommer visas som speciella mappar i din hemmapp.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Sök</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p"><span class="link"><a href="files-browse.html" title="Bläddra bland filer och mappar">Öppna filhanteraren</a></span></p></li>
<li class="steps"><p class="p">Om du vet att filerna du letar efter finns i en viss mapp, gå till den mappen.</p></li>
<li class="steps"><p class="p">Klicka på förstoringsglaset i verktygsraden, eller tryck <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>F</kbd></span></span>.</p></li>
<li class="steps"><p class="p">Skriv ett eller flera ord som du vet är en del av filnamnet. Om du till exempel döper alla dina kvittenser med ordet "Kvittens", skriv <span class="input">kvittens</span>. Tryck <span class="key"><kbd>Retur</kbd></span>. Ord matchas oavsett skiftläge.</p></li>
<li class="steps">
<p class="p">Du kan förfina dina sökresultat genom plats och filtyp.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Klicka på <span class="gui">Hem</span> för att begränsa sökningen till din <span class="file">Hemmapp</span>, eller <span class="gui">Alla filer</span> för att söka överallt.</p></li>
<li class="list"><p class="p">Klicka på <span class="key"><kbd>+</kbd></span> och välj en <span class="gui">filtyp</span> från den utfällbara listan för att förfina sökresultaten baserat på filtyp. Klicka på <span class="key"><kbd>x</kbd></span>-knappen för att ta bort alternativet och bredda sökresultaten.</p></li>
</ul></div></div></div>
</li>
<li class="steps"><p class="p">Du kan öppna, kopiera, ta bort, eller på annat sätt arbeta med dina filer från sökresultaten, precis som från andra mappar i filhanteraren.</p></li>
<li class="steps"><p class="p">Klicka på förstoringsglaset i verktygsraden igen för att avsluta sökningen och återgå till mappen.</p></li>
</ol></div>
</div></div>
<p class="p">Om du gör vissa sökningar ofta kan du spara dem för snabb åtkomst vid ett senare tillfälle.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Spara en sökning</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Starta en sökning enligt instruktionerna ovan.</p></li>
<li class="steps"><p class="p">När du är nöjd med sökparametrarna, klicka på ⚙ kugghjulsknappen och välj <span class="gui">Spara sökning som</span>.</p></li>
<li class="steps"><p class="p">Ge sökningen ett namn och klicka på <span class="gui">Spara</span>. Om du vill kan du välja en annan mapp att spara sökningen i. När du bläddrar i den mappen kommer din sökning visas som en orange mapp med ett förstoringsglas över.</p></li>
</ol></div>
</div></div>
<p class="p">För att ta bort sökningsfilen när du är färdig med den, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">ta helt enkelt bort</a></span> sökningen som vilken annan fil som helst. När du tar bort en sparad sökning försvinner inga filer.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
