�PNG

   IHDR    Q   P��  �iCCPICC profile  (�}�=H�@�_S�*UA;��d�NDE�
E�j�VL��Ф!Iqq\~,V\�uup�G''E)�I�E���xw�q�j%��m〪YF"S�U1��N���蓙��IR���>��Ex���?Gw&k2�'�2ݰ�7��7-��>q���9�A$~��������<q�X̷��¬`��S�ጪQ��r9�y��Z���=��Yme��4��"� A��
�(�B�V�	ڏz��D.�\E0r,������ݚ��	7)�_l�c���m�v��?WZ�_�3��W�Z���.����\� O�lȎ�)�r��}S������8} ��U�88F�������=���M�r����Y   bKGD � � �����   	pHYs  .#  .#x�?v   tIME�8zw   tEXtComment Created with GIMPW�    IDATx���{xTա����$3�dB�$!	HH� �(WAD�h��"ZA���=m=Z��s���[m��Vjk,�*��XQ@@�p`�rOHȅܯ3��A��IBH��@~���!�ٳ��kvf�o��6nDDDDD�W1�
DDDDDDDDDD��R�Hof�����ooo�V+f�Α�T.����z���������:U���E0�1"�������Pe\媪���ˣ��J�!"�  "r�=����(BCCUט��"rssq���&"�  "Ҍ�baРA�
p���$==�ө�� u��^�d2)�����c2�T""
""��K�����Q�����Wcz���P|}}U""
"қEFF�z�~���DDڡ���5�n�w�KP\\>� C�!""�C���㏟�5w�}���3gμ��Ο?��S�2h� ���!;;��kײq�F�e���X�hC���ˋ��L>��6l� ����s���_������Z��q��r�-FC��ѣ�\��tj������l�π������F�~�������ϧ�������C�e�ҥWu=�y����QSSCII	0b����x�� �4i/��"f����Zjjj2dO>�$!!!�Z�
///&L� ��c�:����I�&�r�HII�O�>\w�u$%%��O��7�t��/,,��������63@��o�a޼yTUU�������{������o4�/$))�|���X|}})//'++���{�����Xn�ܹ�~��4��Lzz:��_|����{F�ɱc���ϸ�{%33�W_}�Cgҷo���/�Ljj*n���c����/p��7����L^^�<������׿f	<����[���y�;����h&M�����믿����'x���;���DDD�7�Z��~Meee��}��'����?��?�<yr�^���ǯ�k�v;�N�"77����F||�{�1��^ <���d̘1<��3������z�wȐ!���q��!�v;qqq������~��ӧ�-�_��W��)))���c�Z�����&::�������ƍ�0a��ތ;�M�61o�< ���;�~��_�ּ����Y, @DD���R��k@S��+,\��o����~��;wv8������/�@ZZ 6��>}� �=���ʕ+y��7X�l���wy衇��㏩���X��e���ˣ�����[X�V��>~���vj���^�V+.��իWejRRRb�\\\l����`�jk����=z��C��p�BF������۷o�N��|�EDDDz�A��裏r��a�x�N�6++��������_�BEE���8p������D���E�X�h��:�v;4����䐗�g4���󉊊"66�S���;��F~��_�q�ߤ�|?_���n7?���y衇�4i$;;��;w]�:; ��nJ""�  "�@CC��^������MBB�~����m�駟���g򛫯�gٲe,X���ÇɈ#1b#G���?����[�n%''��zΞ=���������۷/�?�<Æ����g�}������g⃃���CBB��

�ӧ�hV�^�ʕ+;���}j;��駟��r������_DDD����� ���ۻ��'v����R�v;>>>!aѢE<��C>��đ#Gp�\��f���X�b������&M����c����$%%q�����:�+�ɓ'/�III<��sq��Q~�_p���errr��Φ��L�<�����TWW3{�l�ѽw�^L&�����:�~���X


��E�_=�f�`�Ν���  "�>��"r�
���F�œO>	������E}}��p}��IOOo�����',X� h�>���deeq��iHJJ��Ϗo���e˖�|�rc�@FF999���1h� 
�����k֠��Z���((( ""��BCC<���e�|�ώ����ѥ����;���'�_�ʘ>���Θ���7�`ժU8����u����Gux�K�.���&''��JTT gΜaٲe��(//O��������5�����A�n��&���:Mee%_|����>��Jii)[�n������k��Fzz:��v�&**���v��Ͷm�Z�733���~��z��Ezz:����C@�/�]��_Qٵk�����b�������f��b���<�����cǎ���Idd$V����|v������7JKK/����銀�\����.�~W���X�d�������P�(��ʬ*�k]nn�*����W%��(�HoVSSCQQ�*�9s���ժ�v�k���;�����k����SUUEZZ��! "r�" "����&==���O�ե���S�N)��t���H���3����"44T�q�9s�yyy
""
""�g�ۉ���O�>���\EEyyy��Ԩ2DDDD:�f����?���X�V�f���\.���444PQQAYYuuu����Q����D�jADDDD������v���HDDDDz+SonQ h��Y��2w~�ֹ�h�7�}W�^�og�����&8�N�>V�V3V��Ť�CDDDD�N���z��N���(-������%M�	
W��D�%��o����ϡ�v��f3��؈����r�{֭�""""r�0��5��f3�///��\deVPTT۬�oj��UZ� 7v����@���������QG������:���Ju�����R[�l�?\Bh���fhb0.Wz�EDDD������b����RΞ��1a�"�#�:x3|D��u
"""""����@CC�Â	�z��=��=>��(ah0uu�8�N��"""""�8�N��j���n�a����_|B .W�B�����H;a��l >!�U{�;t2�[=�����@"""""��Ѐ����>hk�� @��2``����������t@]]���W��R7�6�Y]�DDDDD:��tb��q8�����V?��(�����tRcc#A�v�k|@'�@�@Ч�U7�kVhh�*AD����Ok�����4X�j��v��N�����t�U�vc�Y�% \d@A@DDDD�2����W�^��b��tY����t��dR%��U,����� p�����d2a�۱Z�X,}��������餾�����~�ZDD�'\��zcc#n�???|}}�n��H�L&^^^xyy���Cmm-��f���D�*���3�[�@Sp�\b�Zu��H�C��������s_f
""�f��\.�B���\�Պ��?.�K�!"r5��~��E݁DD�4]p:��xBD��878���G�/""��i�	��^D�*	��MU� �t6�MWDD��  Ӿ�����DD��� ""�>�A@DDDDDDDDDDDA@DDDDD����@DDDbbb���X�~=999��k�������(�����Ho��A"""�,11�aÆ��d����cǎq��!�fiw�q�����ߒ�����gϞe��� �رc	�j�R[[KYY$##8w�I�&��d"33����V�5j������a�Zill��������Ӎ�Z�/++���\�M����HO�+"""�h���L�:���P��멩�!88�I�&1s��V�3y�djjj0�L���2g�,V���s�Iuu5YYYTVVFhh���)S�0|�pl6.����h&O��j[X�V�����ʢ�����p�̙Cttt��kll$22�I�&����tE@DD�����3b� ������p�\̚5���8���8p� ����kL&�֭�����#G2y�d|}}	

��v��u�}ӦM��,v� ___ ���c��� ̛7���H��mݺ���Z�V+6����w܁�f#>>�����������a� n��V����&�(�<III��w���'����:DD��۷�qg�'N�r� 8v�qqq ���{���r
(++3~���Knn.���8.\H]]gϞ%//���(���:?~���'Z����3~�x���[������� c}������
"=\����������Hwk
mihh0~n?�����ڵkٷo999���Θ1c�3gN�u55��N��s̘1


ؼy37n����\�ܺ	Ѳ<"� ��$%%���t������l޼�+V�2D�q����<d��qo,�4�#������b��ݬ_����~�={� �, ����l~ƾ�����`�1�g��?��ӧ�.FMJJJ�@�4X�l63d���"=\�����|�'�x⊗%..�x�!C���Ç�я~�jY���=��Ì3�����rQXXȆx�w�O|f3s��a֬Y������Oee%EEE�߿��>��S�N��3�xPs����Ԑ���ƍY�f��rDD.���
>�ȑ#�߿?��?.���@ZZ�G�������{塞����r�N����̙3 TUUq��QIHH��ϯ� P\\����l63q�D��Ӎ�J�UWWs��10` ����1�L�XQ�1�w����Wz�������ϧ������rv������5�eeeQQQAhh(cƌi7����_���#G�k��	4����h����l\.���#>>���x�����O��s,\��-[�PTTt������q�\�ݻWo��J;v젴��c�В�c��Ψ��#--���P�����򢺺���tv��m,���_�v����#""���<v���1�Oyy97nd	���́=z4����q�\������Mff&����LD���z�E�_{���@rr2��vUUU���[��߿��~��OUU�����ѣG=BB{~��! %%��_���4�N'����9ң�hs?��O8s�qqq��� �3�� ��Op��SQQ�]w�e�g]�`��o��<@vv6&�����3�|��d"''��>��>�����Oʭ��JYYw�}�����|�r\.��{/gΜ��^#11��Ǐ���x�bINN楗^b	<��������/�L^^��;���<������$''_��c���TVV^�u�}��l޼��"W�#G�p�ȑv�Y�vm�'kZv����//�=��ɶm�ضm���7���0�=м�m��JNNf������7�|�q⩤�Do���@���X��*��F^� ���<{�1�Byy9������������9n��&�\?Χ�~���*����R�n�z�oS�Ҧ/���_���o�&M�d���0ֱ|�r��. ���p:�<�e˖1d�^|��6���p뭷�ԩS�/�3f��2x���OR]]��ng�ԩ0���������a�ر��g?�P t�\��o����.$33�'O��;f����LD$22�o����"���		1fڻw/����$��Ցف�k�@{|}}��4������9r$K�,�I�����X,���M!`�̙<��3�r���̝;����{�=��)))F��d2�����|cc#'N��������3{�l�n�JDD�1WvӜ��y�F�������r��SOq�M71{�l��}N�8Ѫ\�N�b߾}\w�u̟?�/�����p���O[��n������?����xbbb�����5k�����̙èQ��Z���j>�FLL�������w�KJJ
Æ��Ǉ�Ǐ���ʍ7�HHH�O�櫯�2.�7����~�o������V+����ر�h�?��������� 0a�ٷo'N��Ǉ�3g�r�ؿ?'O��n�3q�D���q:�������j���o�e���X,>��6�sBB�����m�FQQQ��dʔ)PXXHMM�G�3f����l6***��o�:�P�H�(++������`���ihh 77���Tc���(t���0�/_����طo+V�0�>7o�oٲ��ӧO�x|�M7����>}�x�����������/Wl���M�Gy���B��>�,YBLL�ƍc�Ν���n?~�~���9?t���l�N'���8F�͒%K���@||<������O=�;w�d������s���ӧOn��&L&������C�3dlܸ�hT����Ճ���6� ��~�u�]GRR`��ɘL&JKKٱcG�����ٷop�rw�x�u���:�n2�

��Lpn�wZZ��8p �~�)����v�m����c�*++�={6C�9o��}�!g�ܹ���t�Kv׮]��߿UנY�fQXXȚ5k���̙3���rrrr���nݺ6�!!!������S[[���0���777�3f�����Ç�ׯ�f�2B�ٳgY�nuuu2��ӧ�f�����:��SXX������\3Ӈ�����?��iӦ��닯�/7�p���aaa�^_[! ΝU���{��UUUgyKJJ��;ṿQ֖��L�5z�h�0�w�f�ҥ������ŋs�w���|�;ƌ���_P[[���7ӧO7�6}���<��ѹ�w��Inn. ���7�}��g���n
?M���444�٭���_���ޡ�<�������



��ϧ�����233��^¹�.���E~~~��^HPP�ٳ��i�$�j{mq�\X,��D���TUU��ސ�l6���v���G~~��z��ө����vs��q�N�������욹"�|��6����,[���{�S�kk]MZv��j.��ݻw3u�T���

������X�[*++ٸq#��r!!!������ԩS�\.|||:\��Ʊ�l��Ǉcǎ���ٴi��z+?����Mͻ�=z�ۍ�db���l޼����ٳ�e�<�r��裏x��Ǚ?��/mu�jqqqth�GS��s]�Z>n��j��N�yg���Á�b�;�0~g�X<�*l^��JKK��Y}��!''����v����Kuuu��S���ƒ�����n���DDD�M݁:�\w5j?����+�������������曌7___���?�����ѣ��oڝb��W_%::�#F���Ċ+���m����^zɣk���r n[֯_ϭ��j��o�����t��ӧO��r�]w1a��y��N�10y�ƍ���dÆ,^�ؘ���F��+)66����n=�=�O���1e_��7���T__�f���:q�'N��n�3e�F�EZZ�y�ڪ����c��>}�p��׳a�JKK�s�$t�R������`�����v����H"##���X�V�wV�8w����l۶��ưa�������_��ۖ��j�x�	~�߰�~���q�ݜ={�cǎ�z�j�-[��k���OLL6����<֮]˓O>١}k9H��3�����o�������'88�S�N��?��������6���ٰaC���j������\�ق.FII�qC �VS����y�)--����q������d"00�nHXXf����zp������������tt��Nooo)//7��uC��s�\ػw/ӦM;�s=Urr�y�״������^�v�N'�ׯ7f�i����_��_�e�~��v�w��|��'�AY[wZn�6����ꫯZ=�V���o~�o~��߽��{�fIꈸ�8222���9����p���&Z^9x� &L`ҤI�ٳ��Ǐ��_2a����`�X(++c�������b�ĉ8\.�O�&%%��}����n6o���ɓ>|8���s����΂������ĸ2 "r5���1� �����
�c�L$�;����?Sn���͎�n7uuu��_QQQ����f�)//��Gmu����v�Z��VUU�������f̘��i�7n~~~��/aժU��^��� ��vٻ����^���8���h���KHH�q��������MÜ�3    IDAT�6��C��kkkY�r�5�^/]���y�޽�ٳGA�2��l8���HBCC��ZMWl3339t�uuum���ǇѣG3`� ���q����RRRZMr�ۻ�r������r����ſ�w�\���e�ҥ�^����m���x饗x�'Z�H����+���o� ..�iӦQQQ�G}���Z�=�~��]�:�D.%��<A
�.���Jbb"�|�	eee���y�<&y�s����Ϻu�<^w�ۻ�r�9�kig�j�_L ضm�q���x�����x�7�1c,��W^�M�D��v����$##�cR����l��+Ҳ��Q���dggs��!N�8�q�Ҧiڛ�����o6B@cc#iii�<y���v8̞=���J:��K}���;����D6l0�<�A�u��7�x#������Q\\Ldd�E�eРA6���`�v;N����Z���)))��g���DDD����墢���
ҲkF[�eBCC9r$AAA444����7�|ctA�?�1!B��c�2v�X��U������r���1k�,�rEEE1|�p<x�#G�`6����7=w�ȑ� ǨQ�

����վ^κ]�f���#11��� JKK����-_mm-;w���ѣ�x�뮻�i����0��F#�С<lڴ�����L�:8wu`РAƽw.v{�:���@ee��A�r,��td��󝋈�\�2�@\\�q_��۷�r]��#G2y�d�ߙ�f������'::���t� 0~�xƌ�1>��f����$$$�~��v��O�8�c�3��B\\���|����Lb�q9�5e��P�ԩS��lDFFz�9  ��'����nρ�c�2x��5ļ�λ��c&O���`x�Y����(**:o7�����������ǹ��+̓��n�b_'�����:z�h�����|EDD���������ɓ���]��F�i�|��I>��s6n�Ȏ;8q�D�gЯ��:��z��	6n�Ȗ-[��|}}�3gN����߿?�O������>}�����/7�x#pnJ�]�vy�.''�]�v���
_�rEFFR\\LZZ��T��_=���������4� 7r��v�9x�����އ��JRSS9t��%��f6�	0�>}��,{�q�-��7�i�IG�����.��z�k���o�ɨQ�:��#���y��7uĈ�H�1m�4l6���l۶���f+:v����ϛL&���III�����lڴ�x����}���;[>p���HOO���?7�|����� M�>}���'N�h,WPP�fW��U���>��S�n7�]w��J

��Op�\WR�V+AAAwi�쾖��_�}(--e�ڵ�f��,���ԩS���5�̓��l�h{���濻�]�/����:�kDjj*˗/���c�����
v����o�}��܊��\)���Fה-[�\�)Ϝ9À ���[���������R
���4bz{{{�4h��Ԟ-������ՖW�;f4��^���A��\�~��qW��g�z<w���,sˮ9-g������\�}8x��%� ��ʬY��c��t�q�F
��ؾ��]�r*�P'N����ow��G@DD�����fҤIF������}�v�͛gt����7������֭�����gt[jo����vw�*��,W���ͻ��e����gё}���p�7e`�ܹ�1QSS���ѭ�������������\;����:��@ӌ(���$&&����n7�$�X��뭨���w�%<<���0	$<<�ٌ�ngҤI�[��UC.55��w�흕n��q�ǝ9�}9��^����u�Fv��˹ͧ��0k�,�_\\�g�}vޛ�t��чs�������mݨ��ۻ���58X�#�=)S����\�v;n��̺u�V>�����c��� ��ټ|tt4���TTTx����"22��Fu��%$$x<>s�L���c�7|/W��BG��'�CRR��r�ѸNOOg�ڵ�6��wO��lF���X�A����Ky���o���pTT���z�߯X���K�^��DDD.֐!C�YTZ�I1b�1�d^^���466��Ox߾}�i�].�y�Xl˭�ފ�d"++���J����������Z�甔fΜ	@�>}��;HMM���
��F߾}4h����Z4h��~;������a<������������餾����jc,��*WW��v�>���s���{��������W_��G�2j�(���5kiii�L&���ה����/e{�:��A`ɒ%m ���gɒ%<��s:*DD�8p�q/�����<gffR__�1�Ls�f�2^��rm1�L����wjG��;}���'N� 00И�>88����z��)��(�s��[Άt��)F�����]wp��IS�\��
999DGG_p_�sZ��7���8���mhh�������n�c�Z6l��򕕕|���W1.v{�:��A��[j�0����Ott4}�����ט�������>�j���ݻ���dذaDDD��kjj���"//���l�+	-�ݻ������fgg�����f���ɸ�nbcc���;����\]a�Ν���1b���מ��)**���#))�W������ %%�g1���d"�ݱE�-���rCT�/���n�������O[�iRUUży�tT��\e


��l������mj�K��}����o��"�*�����s97l���_��u���_�l)99YG������
�.�X��ե78w���^�!""""
ע��l~�a�l�BUUUUUl޼��~�cz2�kY�# ""�������������  """"�  """""
"""""�  """""
"""""�  """""
"""""�  """""
"""""�  """""
"""""�  """""
"""""�  """""
"""""�  """""=(��nվ����DD���ө�}����� P__���KVWW�J���@uu�.犈�%q����Ԩ"DD�� `2�hllԇ���\���j1�L���!X,L&��庤+""������
L&�E""�Ӄ@�v�ٛ������MHDD:��vSUUEIII��+""�1^ݖ@�f��_QQAMM>>>�l6}���H�ƿ�餮����j�N'&�	�Ʉ٬[∈\5A�d2��un�.���Mcc#TTT�]�~�4� ///�<�Z�@�0�t:q:��$""���X,Ƹ � ��,4��n��.""ҙ��
��>�EDDDD��FX�����(�������������>��*�y��7ٷo���U���db�ҥ���',Y�Dq��G?b߾}�۷�ժ
����DDD�h���4�{��>�����Cf���7n�<�������QVVFFF�V�⫯�2�[�`.$66��̩S�X�j6l0�y��7IJJ�ȑ#���������	�ԩS���K�ٳ�w�y���x�5�v���/��?�i���r�JF�ɑ#GX�z5�=����|������7S�La�ҥ���p��!^x�rrrZ���9sx��G����(����{��C=DTT��?ǎ���ҥK�Z����+
"""���8^y��v;'N� ;;��}�2b��j�'�x�x �}���t:?~</��!!!�Z��c�			�����~|||HHH��W_宻��ĉѷo_ >���&33����?Ouu5v��Y�fCll,UUU���r�����s������k�����ӧOc6�=ʙ����<�g�}�3g�PQQ�돯ŋ��0��A"""
=Vdd$v��g�y���gѢEL�>��k�����} ���?�����K����e˖�h�v�y����O��?����f��h�"�y�֭[g,����E������������c�=ƴi�8r� �����7���od��� �3��x}�Q,X`tei*�Ŕ�f���/p��73k�,N�<�0�x1?��{�늀��HSWW�J��������ׯ����大��g�V�^��#0�ϝ�\�dI���v��A��p���,�Nff&yyy��ߟ!C��[���Vnn.��� �:u���D >��C �;Ƽy�0�Ls��i�����۷��{����Gdd$C������ �r�p�\:�z�ߜ����H�׿��מ�l����ŋs�]w1r�H���=z4�G�f̘1���?�d2���dee�Z�ٳg={{{���|.f[������~��ֶZgSþ���e9s���Zx���Y�b��������0`��z}!�ݎ������=��#<��c�5
����Çq�\��f���x��W�e����:u*���덎�fܸq�ٳ�	&��' �F:���/��� ��Kѿƌ����;v,���F9�tYDDD�
6R�^����裏��� 77���Fƍ@jj*n����|V�^����},X��#���"<<���X
=f������^�������8w�����S��e�y�


x�wذaC��u)jkky���)((hU΋�oQP���@o��XEE6l`�С$%%a�Z)..�/���^3���o˩S����;���#::���v��Ŗ-[Z�7##��+W�裏�r�8y�$/���1n`��ͬY���3gFXX_|��Em�R\��W�,
���w�u���b�QTVV�h�kRhh(EEE=�,�>��
��5�O����W������%K����p8�z{.�&�4����4}����U@!@�ҹ�n]	P��4F@DDDz��zH� �O�" """"�  """""
"""""�  """""
"""""�  """""
"""""�  """""
"""""�  """""
"""""�  """""
"""""r��T"""=��d�G //�u�����Ͻ�ދ�d�ĉl޼���k���x{{���ڵk),,���//ƍ����������������������[O����Qs[�n��ѣ�v\��n�x�n�;0` �Ǐ'   ��Eyy9�v�"//OA@DDD�_�~���ٳ6���meIII�b�DLL%%%dffPUUu��s��7EQQǏ'**�aÆ�����������vs���qQQQ�����l̞=���zRRR0��������+�CA@DD������b����Hrr2C���ٳvKy�����!C�������ݻwwKY"""��������?����޽{��{���dee���i�����p8X,JJJ8p� N��Wׇ����H�t:IKK#!!���2l6���cҤI��nBCC8}��шs�����@hh�=��dbɒ%��>�����^]'gϞ������(-ZDII	YYY<x���F�~����1��'���OII�*�W�;��R'ͻUWW+d;��]�������Oxx8aaa��_*���H�+++#77���hRSSU!����=""�ł���d2�񼜣�A�,������B`` ��s}�����  ""�C%''���Czz:���S�p�KPnn.QQQ�~��dggE@@ ���dgg��z����?��呛�{E��m��FVV���FW���eJA@DD��***��6���0�MJJ������T����E�3�L�3��wW:TWW���Exx8���t���Ύ;z�{BB�b�-���rC���:�ED�����t�����s9w�_S�]Ow�DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDDDDD���R���t/�O�N߾}q�\���m�62dcƌ�l6S\\̖-[hhh��2͟?���@ JJJ�ꫯ��� $$�3f`�Z)++��/�������3e�bbbp8�\��������/�K���<��S�������iӦ�̙39{�l��'88�g�}�aÆ�t:ٽ{7/��B��QHHӧO7��M�6ۜ?>�{�u�V���4�2e
Ç筷޺"�PO`1��Ž�̀}����'���\�|}}������X�V���پ};�&>>��� ������gΜ9|��'�۷��}�ү_?rss��Lyyy�ٳ��ĠA���� ��[oe߾}l۶���`���OVVV������0|�p:d����+���o��/2d�&M��������f�ʕ,\��իW_�F������KQQ��կx��w�7o`Ϟ=]Z��s�o�>�o������c�޽:t���`���;�Я_?"""�b�P��~vV`j�_�S� �nV]]Mff&.���I^^~~~ RVVFee% YYY���uy���g2�0���\�ӧ~~~������Jlll�� ??���&QQQ����e� ֬Y��ٳ�����OQQQ�(Oqq1[�n��tR__�޽{	���4#M����T��{i2u}��B�������g�Ν��G]�DDDz��BBB��� ���H`` gϞ%66___L&n��K�2�|���)//gݺu ���yt㨬��f�a�Xp:�W�<�!""��������	�j�vKO����j��`�~���wiy:r�̟?���0���Y�~}��gܸq���RSS�  """��l63k�,������4-_}�3f� �]p��] ֭[��l���g����ڵ��Δ�;\��ؗ�<��_|�;v�u��n/O�{9a�F��7�|�-�	#88�ێ�n���Ǯ��H�h�͜9����V����t>��#>��#
�A�W����ȑ#Fw���J�����uuu]~5�|�����DDD�~��QVV�m�&/T���/�@ii)���ﺼ<���8�#.���G�v�{�^y"""�{�������X,|�;�!((HA@DDD���ӧ�t:ٶm[�������ng���:t�K�b�ۍY]L&			��� P^^Nee%�`���:u����rss)((0��,\��/���G��d2���RWWǋ/�xE���6l�q��|/���)--��<x�U�V�z�jV�^�����?��2��$t�����?Sn�2|���\kBCC�Ƞϰ�0��N����n7yyylڴ	�ٳg��w��.-�����o�����Maa!;v�0��CCC�1c6�����.�>�B�:u*��Ϗ��jJJJ����СCy������'==���~�h<>����x���ۗ��bN�8���˻�<#F�୷ޢ������={��/~��;ӧO7����:s��1��3g�x��W�<-=�������bӇ:�ޞ˹s�W~� �n"�;uwP� �^HA@DDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDDDA@DDDDDDDDDD�{y�
DDD�_BB���/q8dff��SOQVV��~�����r��_��={�t[y�v;?��ϙ:u*N����~������R���pV�\i,�����ӧ��w��m�3{�l�,Y@}}=��?�áC���<s�����b����Ƴ�>Kuuu��gʔ)8���[o�Emm��\HHӧO�j�RVVƦM�<����i�k������ ����Ɋ+�?>Ǐ���x�?���r��rK�����'���ۛ�s�r�-����w[y


�z��[ؼys����ˋ_���ۿ�w�}7�V��g?�Y��'22����g,_��;３��l~��./�ɓ'Y�v-������6m{����ߦ���q��uky�{NA@DDD�TTT���lٲ�5k�0{��Y___n��v^z�%���q�\���������̜9�u��u[y�f3.���Μ9�m�4h �}�vȅ�    IDATn��.?�N�>��U�>}����GFF ���<���s��u�$""��"""(((��v���O@@ V����z �x� v����~��.m��W���hJKKY�x1cǎ�������w;v�[�ছn��o�5��U���~�7�|���J�n7�/�򤥥������b��ل����J��󣪪�x\YY��f�b��t:�ap�銀��H73�L�>�����o����� �x�n+��b!""�#G�p�����{����/wk�4�����O������桇�Ga�ܹ�����_���������ϳr�JΞ=���4BCO;�EA@DD�W���'""�h$��׏��2�lwnn.n����*��}F��m�i:۾q�F 6o�Lhh(����V?p��СCٴiS��_#F��n�s��Q >��Sƌ���w����͛Y�h<� �&++�ۂ@ee%��x�p8����� ��)77���f̘���/�s}���Á��޽GWU����s��r�BH�J(��"H� t�����w,u���5횎�Fl�t@�u�v~ߡNk���*b������r��ȍ�$'9�������ᖠ���y>�:k�����ޟs���g�#9͚5+��pz����Q۷o��ɓ%I7�x����#w���zN�={�֬Y#���׫��V999��͕$M�:U���
1k��C�J����5�|�X�"f����y�^H�F��#G��%#���^FB�GXS�r��ziE ���v����O�5r�H-^�XPyy�-Z���&egg����RRR��}�v=��Q�x_�I�����ŋ���*�׫e˖E����G��}�]���hǎ1}�$��;��ܹs%u�gTZZ�z�-[����K꺐��_����o�YÆ���T{{�����G>W��r�����'��P=�m.�K�7U��ؼqƃ   @\ �'�A��A   @"                                                            =��  ���X�e�Q�̱2�
d$gJvW׼�Wf�	��G>�S��Tf��6  �reȑe�]��&YνPB���T���Rp��)|�c����魦�   �lX��~H�k�H��"�� K��e�5��^��פp�6  �?3\Cd��HFjޗ[��*K�]2�Vp�����N���  �߄���d�����3c�l_����|   �~\Cd�y���z�ם䖵�I)!��  ���H�N�ר���À��'%���  �?���+#� ��1Ү�u�7ip�    b���uw����\��  ��Ȉ�.��_�-I������G  ���%w�XX_w��͐aO���?�  ��[�p��M����l͘1C��͒������hԨQ
�B��O�d�uvvƤIZ�|���n�y��a-^�X'N��B�1�x�_>�?}-E�$e�X����?��I���&�'�H}P���C=�D�d�p��gժUr�\
�Ò�'�xB�~�i�^���D-\�PS�NU(�믿��^z)��L�2Eyyyr�\z�W"�W�өo|����v��^�V�\�z$i����$I�PH�6m�����g  �>��C͝;W�;�����~[��Ś3g�\.��͛�z$���D��Ś9s���߯|�H��^-g�zO�����u�S�s.�n@Ơ��>���C���X���Q=���@v�]3g�Tqq�>��è�SVV�����
�ݦ���iŊ�GEE����bV��b�-�ܢ>�@o���v�ڥ)S����g  �>���sN?y�6l�:j
��}�v]}��1�G�jkk#!�j�rc�����)��?{$Is'8k��t��qF�~��E�ݖz�ΏJ����Orr����~������������s�=r�N�ͦ������P=�a�4M�l]]b�ݮ��6�   �_��̙�_��1�e���3f����4��/�Y_��!�xV�6��G�:.*ș��y��%I۶m�/�������NC�USS��͛�n�A---z�t����������zy�ޘ�
��v�Z͙3G�@@�ij���q���   .V�UK�.Ֆ-["gb������M���[�����+�}�vg�Mֈ,�^��Uր��6�����
��J�,X�@w�q���>����?�AL�7���ڷo�x����z�����{zĈ1$�E�Ǐ�{ｧ+V��>ӌ3  �����X�d�555�^�7u�A���;�9sf�j�jU���o��+��$˰i�wŬ���*�����6���[���kcVK]]�$����$iݺur��JK���(�\.��nUTTĴ���L�l6544H��=;;[K|t� @?f�JJJ����t�Ҙד�����4=zT�Es���r{�%GJ��M�:QnWW��n5tǸd�4�����	H�������ږ���O��i/�X���d0@uuur8�5kVL�z766j���<y�6nܨo�Q����x<1}�1BG�9��ݾ��z5`� ������Eyyy�x<�;>]��/*4{��y�#�)E91� @4���ȑ�h[�h�n��f4H'O�ԡC��裏j̘1z�W����|��z�'bROvv��{�94H�pX{��ѳ�>9�|�l_����kz\��<8P��~��;�/+#�OK��d��������
���%o�_��JIIQ8�������F��}�z$)//O�/Vjj��^��-[�ݻwG���o�YÆ���T{{�����G��{�Z�~}�.*�v=#G��ر]w����ڴi������.�˥͛��5H�8�A   .�@��ް@���b���?*���" fb�F   �L��Θmیᶁ��    b���D
v�����
�n� A    &�
��ۡ��},;h   b%�����
x��A�&   �dz�>�����~/�[KÃ @  �X��&�q�C���
�]A�  �/�
n�7���y	z��A���Ag���yu6*��i)���   �7|�
m~JfGϿ���i)�pZ4�e��sKϿLl��+��'2;N�� A   �7��B�5�$���ҭ��~?��LO  @���(��	���~�����-:��7�������	�����U�5Ӯ�C�f/���������Ҋ �+���VCCK	i���_�a3$[b��T�r��Wrw �k.�K�7U��ؼq�#�l�  ���5+����Ю�d|��A��H.9�d�]�$3����d6�Y�K�O��0�    ����m��m�-�K�k    �     �     �     �     �     �     �     �     �     �     �     �     �    ��e�	  ���jڴi���֌3����7s�L=��#�Z�:|��JJJ����Z222TRR�Q�F)
�O>ђ%K���)I*,,�SO=%�˥�G�������Y=j�����Zc�>˗/W^^�$����Z�x�N�8�z���4m�44H�pX���ڸq���`��L��ѣG�W^�j��TϷ��-9��)IZ�n������{�3  �~���Ν����nӇ��{L�>����N;vL�<�HTk1Co������5g��\.͛7/2�'?���/_�Y�f�����?~L�9_�Ţ��j�E�������X3g������`���׳o�>�X�Bo���ƍ�m���+!!A�P�O^���y�w�b�
�X�"nB A  �~���?WCC�Y�

TQQ���:IҦM�T\\�ZN�<�6(
���k�����ʒ$���(++K�ׯ�$�\�R��zk��P�Ţ��j�E����F:�V�5����ޮ�G�*+
���F.�+2�f�iҤIںuk��^=��  �c�V~~����d�n��Veff�b�?��Cs���ڵk%I��٪�������Qjj�GLꉵ��ZϷ��˗k�ƍ�2e�^x�>��j�jĈ*//�L�0a�����ggpz�G�fϞ�{�WEEE���  {uuuZ�x�/^��_~Y���
�B��x�;MK�.Ֆ-[�a�I]G�c�\��҅�E������}M�6M[�nՃ>�7�L�E_���t��q=zT�������<x��;��G����?�7�ЪU�����I�&  @��n�:=��Ú;w���٣��ʨ�Ţ%K������䚚eggG������x���cRO�:P�'��f��`P��fΜ�z�������ѡm۶E�ggg+##C�����~Y�V��������cR�$���H��~������\�	w ��:t��?���t͟?_+V��z����D>�OK�.�6���Juuu�>}�֮]���[k֬�Y=�p�zbQ녶������4=zT�Es��QYYY�k�6m�B��6n��m��]��k׮��y��Z�*�w�P=v�]�Cmmm�aC'O�����Pa/)�g<R�#���74 ���v���"�E���o֠A�t��I:tH�>��$iٲe?~����s_|�Ũ�3f�^y�544(K�>��S=�����#Gj���0`���˵h�"555Ŭ��]_��S�}]Ovv��{�ȭ3��٣g�}6r�y4dff�������#����j�[��ey��X�"�A�B��\.͜93r�KMM�6o�,���'�{�˥͛��5H�8�A   .� ��� �5   @"                                �}0h9    ���!ɤ�   ��
�     � Â   �8�    �0    �� �Y     � �    q    �Y�l    �A L+   �8#    �a    @    @    p�~@   �� ��   @�B    p���=�aA  �������hԨQ
�B��O�d�uvvJ��p�BM�:U�PH����^z饘ԓ����_~9�lRR�jkku�=�Ĭ}n��V}�{ߓ$��~=��3ڽ{w��9s�y�Y�V>|X%%%joo��{h�����˓$>|X�/։'$I���zꩧ�r�t��Q=����x<Q�'99Y����Z����Tyy����$)77Wiiir8ڹsgdz,��l���Wrr�$���E���
���w��X �3Co������5g��\.͛7/2�?���v�fΜ���b}��1����N��őǺu�bZ��f�SO=������7���^{M�=�X��2d�{�1=�裺��;u��1=��#Q������X3g������`��ȼ���'Z�|�f͚��j���Q�'//O���ڽ{����5dȐȼ��&�߿�O;���0���k���ڽ{��V�����滇   @��<yR6lP(������ە��%��H�wܡ�{N~�_�pXUUU1��t����1c��{ｘ�c�X����i������SPP���
���I�6mڤ��⨿�jkk#[���������,�_�^��r�J�z�Q�%!!A�C��͒������G�{�^�>�|]��@  ��#�4e���^�G�|���� ��p8�3g�~��_J�����&͛7O7�p�ZZZ��/���1��t�7����H�7���~-Z�H���o��ze�f��)}]��Ç������<UVV��[oUfff$�D����5f�UUUE��ggg���N��5����F���r8���Qk������e��dF����L���Ţ�F=h�'���"a  b�j�j�ҥڲe�6l������}���Лo���>f��n���Z�zuL��n��;�������j�̙����/-]�4f����i���Z�x�^~�e577+
�I������M���[��������z�0���%��O�� �E�  ���Ţ%K����I/��Bd������%I�֭���VZZZL�9%;;[#G��ڵkc�>cƌQbb����/Iz���5~�x�����Ϻu����k�ܹڳg�*++��Hx0�;Ｃ�3gJ�:���	������ �����k���`L����S! ��������W/  �e�JJJ����:���ب�۷k��ɒ�o�Q���Q=jy�zN�={�֬Y#�������UNN�rss%IS�NUeeeTǠ��>C��$���k���Z�bET�'555r� �Ţ9s樬�L�TUU���:M�>]�t��wk͚5Q�������G��A������WO����)���2�{T��xf��kJQ��^/�� �+���VCCCԷ3f����+jhh��#���O��OD:*�/Vjj��^��-[��c�T�$���*))ю;b�>w�y��Ν+��B�g�yF���1�gٲe?~����s_|�Ũ����s�=�A�)kϞ=z��g#g�F��ŋk��*//עE���1���C��򔚚*�ݮ@ ���:t(&�8�N�9�[plmmUyyy�|Ǹ\.m�T��c���>	#��"   p��    �k    �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �    @    @    @    @    @    @    @    @    [6�  ��8p��O�.��!�ǣ�>�H�����Y�f)--M���ب�?�Xmmm1�產�"�=Z/���Y����{�G�C�iJ�֮]�����c��4e����+k���ڱcGL�q:����;#���v���j�ʕQ�'99Y����Z����Tyy����$)==]��$�����ʨ��/TOFFF����UTT(  @߸�[�}�v���kҤI�0a�6m�$IZ�~��^�$i�ĉ�8q�֭[�z$i���JHHP(�y�HҪU��ޙ�m=7�t��V�^{�5��a0 f������^�\KKK�����Suu��������!C����R�a(??_{����SFF�rss������p8����}�����+''G�VUUU\|�04 �KII���Tyy�$i�޽�ꪫ"�O� �0d�Xb^��f�M7ݤ-[����O���nWaa��l٢P($�4����m��l6����Q�'!!A�C��͒������w�����j�*Ĭ���$uvv���K�<�222�滇3  Ę���v4���*!!AV�5r�}֬Y���RKK��{ｘ�s�7j�޽����7�3g�I���ǵm۶�v./TOJJ�:;;5~�x2D>�O[�n�ɓ'c�>�4|�p���G�e�8�H�Z��~�l6�Ði�*//Waaa��Ĭ���%&&*11Q�����Ȑ�n'  ��q��t!���,�&M���c�j۶m1�'33S���ںuk�i�?��jii���дi�t�M7i�ƍ1��b���r���A[�nUAA�����bŊ��$���0�CpzSkvv�<���v��nD=�����ѣG���/��@<ah  1��z��#w�\��|g����ڷo������3x�`8P<��x�Y�V�u�]g����95�������TYYY1k�SG����$I���JNNVbbbL�?.�Kn�;2|(ڝk������P0�i�r:��X,joo��u���a1�G������~�߿_���Q��    "ZZZ��zUPP I=z��9"IJLLTjj��������jll�Y=;w�ԫ���+VhŊ
�Bz������z�v��N�����#F�PCCC�ڧ��C555:t�$)''G���Q�\^��S
u�ȑȝr�������G�t5hР�����+!!A			����T�|�^�шF=�"��l62D'N�����Pa/[�<�֔����3  V�nw�;��ok���JHHPSSS���.�K��v����e��N�8�-[�D�����9�������^��Q����߮�������jm޼Y>�/f퓖��[n�E������ڼy����b�z�{�Z�~�jkk���|��u����Y�P(�cǎ����Ç���$��׫���Ͼc\.�6o�Rױy�A  �� �O�� C�   �8D                                               ���    IDAT     �$M    �Q �Yu���   �x	 �L�����N#    W2�b��h��=�f���o0�i   �+7 <��"�q�|�    p% �ФI����)��ꬳ�2�׿�   �+����4�;S5bD�9���Q��ŏUv��     \�F��o�+ҵ��7 ���:t�62�     \�F�����.�ر��9���J�}i�v�:v�<�    p���W����'kҤ�� ���Y;v=�:   �e�`� �w�dM�Zx����W�w�w��m+�q]   �����������!�������mզ�e�f��I    ���au�7�#e�XΚ��I����
    ����J�=�ݤۊǜ3 T;�7����~�O�p�m�   @�]�Q: �'�0��:e������n#��� PWע7^ߦ��� �   } B���Pbb���V�%�0 ���;
)���C�i�j�~�@0��ҝ7Q;k��g�?Qߢ�WlӇ�V(�$�@   J��`0(�4�t:���L� W�0d��d�ٔ���������b��n��z=$��Y�5���r&E��)�z��O���T����@   J! +--M��F�pII]������
�>w�\�$9�ݻ�O��^��~��g��Q��   @��a�\.B G�\.����E<���Vo����]z{�'�h�G�^�   �Щq�V���@@r:��x<���N�V�ީU+?Q[��Oj%  p��B!�\.@�:}}�A���z���|���y  �옦ɐ  ���>��Z<�} N���  \zg�� Υ���m  �~' @G                        .��  ����I�֯_���: A  ����ɓ5l�0I��ի���A� ��   q�3  �cV�U�ƍӰa�d�����9���Pyyyr:����
��x<:p���?�m}cǎU^^��PUU����u�7Jb�@   �����u�UWI�|>����5dȐ��8p�����&��-�ۭ�?�X���g����S�����ɡ��   �/���4|�pI҉'���K��M�����n�n߾]>�Ov�]�CV�U3f�PBB����T[[�m}���ڰa��8��   @�����0IREE���$��ѣgu��1c���t�������WYY)�4e��*** A   �G�iF�}*�2`� M�8Q�a���Aeee
���������o}��@��A  �S�'�I��ʊL?��R�#�������PCC��v�yח��+�0d�XTPP@cq�3  �S*//���Õ�����$I:kOss�B���V����:��n����b������2]}��2d��̙#�0d�Zil qF  �~��>SYY����p8��;wv[���j�֭�x<JIIQ^^�8 ��{��v�ءC�����f����N�w���B4:'C��h��kJQ�9�d  ���n544\�sLӔ��;k�N����`0�@ �?CEEE2d�B���}���< _�����r.�K�7U��ؼq�#� @���Ԅ	��ب@ ����ȝ����K �A  �8��z��Ԥ��T9��թ��Lǎ�� �   ��<yRk׮�! p�0   @    @    @    @    @    @    @    @    @    @    @    @    @   _����=�Z�J�֭��w�M� q�F  �?<�裺�[��o~32-==]O?������p�B���\�m�;V��{����I�����|� @��   �Tnn���?�C~�_����x�B�$:T���ڽ{��^���Z���1E�rŧ �~h̘1Z�d��o߮��~:�Q�X,��������r�ݪ����ի����N�iJ��|�I��a=zT��~��N�v�ڥ�^���3fH�֭['I�뮻��ب�n�M��ַ������FmڴI���o���Y�$UWW��[oUFF�fΜ)��߫�^�.I���k���}OÇ��bQmm�^z�%mذ�7p�qF  �~f�ԩz����?�Q?��O����{����W_ռy����k޼y�뮻�����H�PH=����^0@,�$���?���s���h���>}�u�wj���z�����o[��o��1c�����)S��4M͝;W�f�R ��s/T��f��O?���R}���ռy�|�ry�^�@pF  �~$==]%%%z��7�|��n���<�7�|S���$��������C=��+WF�=~��^{�5I���׻ﾫ����ݮ�bѷ��m��W�Қ5k$u�����_�J���jjj�$�8qB�����/�����r��t������%I����) �   W���V������o����u���ȼA�E�Ӝn׮]����5p�@�<yR�TYY�m���&%''+11Q���gmw���JIIя~�#��G?:k~NNN�3_^^	�����ܬ?��OZ�l�v�ء�;wj˖-:r�o�   ��-�_��_���X�?���q�ܹSR�I�k�t��P(t�eN��LK�h����k<�C�ܞ�Z�l��z�-M�0A7�p��͛�_|Qo��o��  ��@ �'�|R6lвe�t�M7I����֦�c�v[���SKK���6�����ڪ)S���s��ȑ#z��7�p�B����={6o
 
8#  @?������jkk�O�S=���Z�v�V�X��s窶�V�w�����u��w��_�R��B��o�G}T�G�ׯW аa�4u�T=���Qy��rssU\\�-[����N���7n����yC   �i���/)�׫E�)99Y����d�Z�����v�ĉz饗���o��Z�J�����7��{�G�`P555ڸqcT�{Jgg������JMMUKK�>�����'o 
C�f/���x�5�(�[z �Xn�;r����|>eeeр@��x<�Z��ri�*u��7�xD�    q�                     \��  ��#F���@���*++����/j���v�&L��!C�(���Teee���}���땓����D�������:p�@���    �T{{�v�ޭ��܋�o����F�A�7N���z�������S����E�������h�ñc�t��0@EEE�x<����7� �� �O?~\���
=�f�i���r�\�X,6l����#�ϧ��zUVV*??������jkk�����U0����W� ��  p��裏���*��)�ͦ�������f���IR���������p8��zu�ر�n �   �L�TCCC�w�-ұ>%�n��j~��۷O����VFFF���i �   �wNu�m6[d���n�����g�={�9����B�UVV*33S���ڻwoT� A  �+��j��ѣu��!���)*555r�=--M�G�z��:��a���Ng���ٸX �~�0Y�VY,Y,Y�V�ѫ��E�\s����*++5z�h98P���������Gk�v�F�!�ө��:T���:q�D�� ~�sTh�2���kJQ��^/� �"�������2MS>�OYYY��k��V�F��6m߾}ڵkW��.V��P�V�UEEEJOO��fS[[�>�C��s]�� .W�=3�r��yS����g<  �M @�� ��         �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �   ���j�ҥ=N�޲�  ��>�����^�Z{��QRR��   �����I�=�X�i�G���4 �   W�P(�Ç�5}�JMM��?~��>��
�B:x���n�\.m޼Y?���4q�D}�;�QVV�JKK��3Ϩ���  �J0q�D�A-Z�HZ�h��z�)9��g?S8ֿ�˿h��*))�� �   ��n�֭[�m�}����緶�jٲe
�Ò�?��Ϻ�;t��w���I��r�J��?��  @q�kN�<���>|8$���A�pjZrr����I�  k�F���@�����`0x�4I2���#        �I0i    ��
{��3aM)ʑ�� W$��}���7MS>�OYYY4 �<O��s�\ڼ�J]�t�3���         �     �     �     �    �˔�&   ��V�Ǝ���+))I���ڳg����"���vM�0AC�Q Pii����ι�����u]�}��>�z����1�~�=�԰a)����" ����������~^(��庨��l6eeeiϞ=*--U(�ĉUYY�[{�7(99Y}�����5i�$544���]�a(33S>�O�p������/��}�i~��R��|�Z��p�Xe���~G  ����g����Q���:|����ڔ�����bѰaôg��|>��׫��R����N�����r�z\����ڇ����} �	A  �~(11QN�S��͒$��)����$577+55U���G�����e{��}�i~��J�5  �3�E�'OVYY�ZZZ��`�l���)�@@v�]�d��z�lO�=��o� �q0$��  }��կ������?�L?���l
��.�=������ŬK�fϞ}����.jz;?� ࢂ !  ��d�&O�,�0�m�6����-nkkS0Tjjj�yZZ�<���;�=Z��qٞ���������h��s�v�  ��n��&9m۶M�a�j��0���UYY�ѣG��ph������UEEE�t�E�\s�G���4?Z������@|}侮����3aM)ʑ�� W$��9��[�i���)++뢞�t:5k֬�����:x���;=�Co�1�� \
�=3�r��yS�������C	  �  � ��                                �g��E]    B�� �   @����4 �   񦽽��A@��>�  .1�0���Ac q�r��  �ĬV��PKK�|>�	�ϧ���   ��0�H����F���1L�������v555]Vu�x�  ��,K����ڪ��%%%)!!�[P p�v�C��|>����#w
��>�  .1�0d�u����2MS�`P���jmm���+�so�,��g�A  �(��P(�P(�� �
��[�VY��˪n�   Q�H�,; ��g�    .�����]�    �     �     �     �     �     �     �     �    �◅ �2�4i \n�"N   � 
�0%&&��p�j�^v g�C����:::d���V�e  D��e���N����i�
b�l6�l6������ѡ��VY,����b�F  �(��p8���TB �������P(t��L   
��\.���	��!��E   �7l�Z9 �!��I   ^�B!%%%�   ��4�   @<:uA    G��                          ���&  �򔙙��ӧ��>�$]��Z�n�N�8��s������v���I~��y����QQQ�$i�������Um�]o�����~�    ��iӦ);;[�PH�W�����6ʔ):t�L����utt��󩦦F^�W�TSS#��Gc   p�(++Svv��V����t�Сȼ��2D�T]]���I���ц"������~���;զ�i�   ��S]]���N%&&����[��ϗ��uYߑ#G$I�����˓���nW0���сt��qI݇�:tH�F����<��ժq��iذa2C����
����ѣG+--M6�M~�_���:p�����λ"egg+hӦM��d������J)))�$�׫��r<x�[�;??_W]u�RSSe�Z��ޮ#G�h߾}UGo�y�6mnn捌�
 ���aUTTH���ӕ���WPP Ijoo��8p��UUU%��'�ۭ)S�(;;�ۺSRR4q�DY�V���0~�x]}��r8
���������-c��u��7+33S���V{{�222����c����k�����aܸq�0a��������������q��i�ĉ�宻�:M�4In�[�a���U�C���]Go�y�m
�g�  ��8r�F���755i���JMM��?udz�����|���r8�Z��1c��������n�O?�Teee2�Ã���4|�pI҉'���K�v�������}ضm[�(��j���`绣�C�ׯWKK�y���t�k��$���F�>M�4Iyyy���������#m��Ԥ�������0�s����m655]T�  �+������נA������;w*??_R������Ȳ�֘1c�t:�ZOrrr��wvv���,��s�eOMM�tf+**�%IG��Z[[��ޮ��d�v�m���jiiщ't����֛������B!�]�6ra��dddD�8z�h�֊�
���E���|��N�S�wz��7u�v����7m
�w �9չt8��ˋtDkjj���.I0`�&N�(�ө����/��͛���)���O]\�[�wjO�SB��֬Y���R��������vkԨQ��W�zֺ���LӔ�j�W��Kv��b�s���6  ���;��q�d��%��E�R���������PCCCd�/���D@VVVd����$��&�ͦ={���?���kϞ=�����V�رC�4|�p]������1RG^^^d�ͩ3#��9}�k��F			��p��A�����4 �	��:z��F���wvv���:�Lss�B���V����:��n���F�,�Ettt���\ÇW~~����$�ot����Ummm
�B�eN�P��������3f����j��a}���笣��M�҈#����ٳg�4��p����������+_��2224k�,y�^%%%���)r�Co긘mW�  �ϜtJyyy�����֭[��x������<8p����=���TVV�@ ��*k�Νݖ����q��܆���\[�l9�KKK��~I҈#4v���.�c�m߾]MMMr8JLL����Ν;�׿�5�ܮ]�����E2MSP ����WGo�	\IC�����<�֔��/�� @�v����pQ�1MS>��!5 �����r.�K�7U��ؼq�#�8#    �!�    @    @    @    @    @    @    @    @    @    @    @   }c�Z�t)�M  @�������O3f�Pff�:;;USS�͛7��W_���z��Ǖ������ݦ�ٳGIII�q�ꫯ�ܹsu�5�(;;;�^X�`A����oi����\���s�^�ZN�S?��O$Ik׮�|�Y�f���HJKKSGG��;�w�}Wk֬����p�;��m�ݦ��K���߯W_}U;v�z;L�:5�]I
Z�jA   D�?��?k�ĉ��ٻ�訪���ߪJU�"!d 	C ��y8`#�j��B��m�[�.,��4������*
/ �ī�2#  Cd �ȜJ���Gn�KH ��V�U�3>����眽��;w.��f�Obb�uۇ�+W�@4Am۶eРAdgg�t:������>���]�3��SQ���_�~ <x��￟��gϞ%::���P�u�FXX�}� /��"����g��5kF�>}�ի3f�`�֭u^?��iiiF����z�d21x�`,X��ի��8P�r~��73f����Z������GU� ���x�^��Ҹ�{fϞ=��_�����<��:�u���}5wڴi���2cƌjo��Ϗ?��6���֭[ٽ{7�'O��;��l63f���^"""���e���,^���W��m۶1b�JJJ�?>m�$��    IDATڴ����w�fʔ)�^����3g������ѧO^�u ��.>��3Z�n���X�d	���`�ܹ$%%1iҤ�x�^#�i�����>��3g�гgO���K
/:��ngŊ�����z2d�f�b�ĉ?~ܘoРA=z�q��a�٘={6O>�$/�����6��M��f{�ƍc������<x��裏VY�o~�Ǝ��o�͞={�ݻ7�'O��v�t�R� 7Xqqq���ܹ3�V�������ɗ_~ɚ5k�z�2b� �����㏫,�g���˱�lƶM&S��2��|ߦM���9y�d��E����޽;����۷���%"""R�fϞ��������9z�(`���lܸ�����J�1�{��;���?4>�����O?5*c_~�e���V����f3�G�f���|��� |��$%%wL&cǎeɒ%�Z��ؿ��hƍ�D�r8���MRRS�N%>>�w�y��w�����f���zY�h�qN���ЩS'F�MϞ=���U��GFF�i"p����V�Zq�m���7�PPP�D@DDD��޽{���~G��ҥ]�ve�̙<x������\.���y�G�ѣaaaX,���9u�T�u���W�;//��� (++��>]i{����o߾*��߿�H"##��I�ڳgcƌ!<<�3g��h 6o��?�`���X�|�M"""x���裏())���V��I�&1j�(�n7��������1}�t{�1@\\l޼�h2t~��k���@߾}���e�ڵdee�����M�6JDDD���|>>��Ç���/�ꫯx��72dk֬���;�����:u
��ɴiӌ��.������Q��]N�6/�@}����*gee�c����b!""����ŋX�p�1�Udd$/���;w&//��^z�ݻwWY_~~>s�̩����Ӂ����o�Z������z��cc������c�W(�7oNHH���̟?�]�v���M~~�;v^����b�\v��l/77���R�v�Ze�.]��srr())�gϞU��ѣ����={V���0a			�߱���t�M�9�����d"  ��� �V+ �z�b޼yt�ܙ����� ��Jo�ۍ����ot8߼ys��2Ԅ�b!..���@cĮ��h�������z�>��o��ȑ#�={��-[2v�X\.[�l������|���Ǯ]�0��L�8���(8P�㦛n"..���|�ѱ�Ru���zY�t)����8y�$�b��8и����X�`�Ǐ��ɓ���/��ݛѣG�������=z�`ڴi DEE���Ȃ �9s&ǎc���<�裔��PPP@tt4fs�u�E�QZZ��n7�����0e����gT���<{��2d=�������k$�o��V����d"!!��n�	��DQQ[�li��֔�����֭#99�Gy���`


ؿ?O=��1��/���ɓY�l�����6�x[+V��{����;Ç����Vk{�|�	���<��3��.d	�<�/�b�0a�"""�����?dٲe:��@@@�Q�d�ٌ�l6 ���g���$$$I~~>���|�����F�~�ĉT����y��*�p��a��Ӊ���f����ͦM�X�`��T����ڵk��q7�H�f�'�y//ɃZ��-�)""�ӧO�h�χ��e˖M����еkW�q�H��T�s��ng�T��7���{�# """�$66�=z�{�n�^/������V��cJDDD䚍9�'�|��̉'�3gN�'$��id��������i`4|������Q" """""JDDDDDD�������(%"""""�D@DDDDD��������MӦM����
BD.�OE ""R0z�hn��vZ�j����ĉl޼�e˖Q\\\���ݻ���@�T�}��ǠA�h߾=͛7��p�����_~ɷ�~[e�^�z1n�8:uꄟ�iii|���|��� �����v�Z֬YS���l6F�ŰaÈ�� %%�O>��]�v�y9X�V���Kll,.��}������D@DDD��n�7ޠe˖,X�������i׮��s��%K�Tk]+W��|���ۭB ��~p8�={���hBCC�֭aaa|��g 0�Y�fa6�)++��pбcG�M�Fxx8,��Ϗ~��p������_d���x�^���C�f��ӧ�z�bƌlݺ��c�����ϏC�]0�W�^��W_­��Jaa!���JDDD����O�u�����ĉ��G���o��y�� �|�͌3���x�V+iii|��GU*IӦM#44�3f,���,�J�->|8n��1c�p��Ann.˗/g����|>�&b���̙3��������ӧ���: w�u�QQ�4if����,�qJKK�={6���c	�\���Mu�ߺuk��%K�7o s��%))�I�&�J"��߅U`��L۶m���q:���撞�N�v����H�C����;�d͚5U��s���wV�XAjj*^��!C�0k�,&N�����/����d�,Y����p�\����e�ر�����ٳ�޽{3y�d�n7K�.Ձi">���*�ٳ���rl6���u�ִn��M�6��������J�>}X�n#F� ������7�LU������mڴ!::��'O�I���g|�*�sqqq��wG����ȍE@@ ǎ���֭��׻wo��>���K.��������z���رcY�d	�V� 33���hƍ�D�	{�ᇱ�lx�^-Z@˖-��gϞ5ޟ9s�x߲eK|>���\l�������ЩS'F�MϞ=���F_���ȫJ������2���D��X~��#�8�ɜ���j�*��!<<�Gy�=z��b!88�S�N]v�cǎI@e�*88�={�T�oϞ=�3����*�<i��V+�&MbԨQ��n^y��9ιW��e6�ke�>���ӧ��c�1`� ������`���F����ײ}�vc?;v��b!%%��NT������e�o�{%"""R'rss)++�}��W����;�����:u
��ɴi�.���\N���ߕ�K�P��%22��^z�Ν;����K/���ݻ���^�oѢE�ĴҩS�		a��� ,\��O>��Z뇊�8s�̩����Ӎ
{FF�U�v��r���|8�*󔔔�v�	���� 4oޜ���F{���z��r��w�q��wӪU���ӼysBBBHLLd����ڵ���l���iӦM�����CII	={���y�=(,,���C�^�z1o�<:w�LJJ
�?������L�"~�-�`��1���y��9�s�NL&�j��~����v��w�����o޼����^��Kzz:]�v�f�N�6m.�說��z��ޣk׮̝;�p��JJJ��C�l��ҥK��ϧ_�~�ڵ���ĉ������5ڞ��c���?��'O��/�лwoF���￯҄L�2���0 :t����i���<��� ���̚5���X>��3�N'���@E_���|�v�1�~^^^��?d�z�!233���'66��c��[o�y9�ڵ��}�2b�\.�w�n�#)�G
y�'x衇�կ~ţ�>���"33�����+W��zy��<y2˖-��p���߳aÆ����ŋ�X,L�0���rrr���Y�l�Hr�{*�l6���-[x��g��q��>��sV�^mT�'N�xU�?|�0������`�����fӦM,X��H*���f����͛��q'�� }罼$jU��hDDDn�����pu�|>�Ng�VD�i�n�����'�h�o:�U��G@DDDD�	R" """"�D@DDDDD�������Q" """""JDDDDDD�������(%"""""�D@DDDDD���������_|����o*�1?���H�0i�$n��vz�z�?3f� 00P�FѫW/ƍG�N����#--��?�����ژ�C��?��;�޽{y��'�y���y���X�v-k֬���cРA�oߞ�͛�p8�����/���o�5���l�5�aÆ@JJ
�|�	�v��2���[���\.>��s%"""�4����v�UMȀ�5kf����2;vdڴi����`� ڶmˠA������t�����_�~ <x��￟��gϞ%::���P�u�FXX�}�Pq�k���x�^���C�f��ӧ�z�bƌlݺ��c�����ϏC�]t�O?�DZZ >��q�uꋈ��O7�|3cƌ!>>��JZZ}��e+C111����رc̚5��={^q/��" YYY:�-Z��7�0t�P ֭[��9sX�|�U��o�&M�l6�����?Nii)�gϦ_�~L�0��+W���϶m�1b%%%̟?�6m�Tk��ׯgΜ9�߿��G�>}x����뮻���hݺ5`ɒ%̛7��s璔�ĤI�j��������U`�׋��iI�N}���n��b�
RSS�z�2�Y�f1q�D�?~��III̞=�������^����HNNfɒ%�?���2,�E��t��~kݺ5�[�`ӦM���ү_?�V+}��a�ڵƴ�),,dĈ ������W�gϞ=���c�ٌu�L���������l6޷iӆ��hN�<Y��ѽ{w�w�Nqq1���#''G�����\_�W�+}�����ݛ;?��ʴ�2s�L>��#��EM֑�������zku���kٲ����ٳ��3g�\t�+��|WL~�al6^��E����IJJ
�:ub��������^��~dd�U%���DEEɅ�d�C�F�?�� G���p��xhժ��v�|�JDDD��	�G�G����a�X�ԩSU��ѣ��~;���
k֬��u;v�ZI@M�)ùW��e6����V��I�&1j�(�n7��������1}�t{�1@\\l޼�h2t�}W�o�n�ӱcG,))) U����,�}aa!�i�F�����\_���)--��w��ԩS8�N�M�vA�挌���������q85^���������+�-Z����U�I���ŋX�p!�|�	Pq5���^�s�������K/�{��*����3gΜ*�M�>ݨ�gdd\U���.���W�{r)�����# ""R����������ٵk������_�sf^^O?�4AAA���k�����b�n7���K���L��}�-�`��1���y�F�y�Ν�^��d"  ��� �V+P14�y��ܹ3)))<���$ 			��пc?6o�\�>
W�b�G`` 6����x������n��^����H=T\\L~~>���c׮]��f&N�HTT�`���B�y�������{������|YYY�t�M��ő������~I����2k�,bcc���p:����}@���fhӦM0��'&&ËΜ9���\RSS�$`ʔ)����"����\��2d=�������@nn.o��V����d"!!��n�	��DQQ[�l��WB������	��b[��zy��<y2˖-��p���߳aÆK._RR�s�=ǬY�x�7x��gk��s�X���ݻ��;�lz-��i˖-<���ł��8r���9�W�6�0*�l6��Y�(@'N���mT>�kBf�ٌ��&==���l6���lڴ�Iŵ�T��v�Y�vm�:�&I�l��;��%yP�:�E#""r#EDDp���-���p:�5e���/�L�-�<y�
_��n�b����'�h�o:�U��G@DD�kӦÇ���l۶M""ׅ�����`�=�����^��%K��@DD����HS��E� "ם������(%"""""�D@DDDDD�����%�|>��(ij*�,"�D@DD�	)//W!�������T̓D�����W" ""R�L&n��á�ib��^����H-�X,�L&
q:�*�&��tRXX�D@DD�)2�LF" p��YJJJ�LH���|������נ��O�NDD����f��_TT��� 00�*���4�ʿ����tRZZj�֐��JDDDj��d�ϯ�_�������v�)**���H$�H��&�	���4�Q" ""R�ɀ�����y�H#��[,,K��o%"""uX9 dAD��;�D@DDDd�@D��$""""�D@DDDDD�������Q" """""JDDDDDD�������(%"""""r���"""u���D����q%"""u� x<L&�l6,K��0�ȅ�o�ǃ����p����X,*!P" ""RG��ۍ��#88��� �H#b2������Ϗ��@EEE��f�Vk��A}DDD�(	�z����*	ii޼9�����:��z����l6�Ha�ٰ��JDDD���v��EwD����`%"""M���!00P!"JDDD��ϧ&A"�D@DD�)�FPDD����H����Q" """""JDDDDDD�������(%"""""R;�T"""STTw�q;w��O�>�[�����K.ӪU+���ϩS�T�Ҡ��׏�� ~���k^W���i޼9k֬a���9s�m۶)��s�m����a��唗�W����L�֭��|�X��Á��$;;���b ���q:�*L��z��Mbb"gϞ�����[e��n�{��d2���r�̙��iiidgg�o�>����1Q" ""R�����b!..�Ç������� ++��@AAA��������i>�OQ������͛F^^��yBB������'O�4ާ��7��D@DD���ʢ����� ڷo_%h׮fsE���G����D\\���X�V�n7<x���L ,�z��m۶�L&���.��]�vt�Ё��PL&���<x���4c�;３�����8|�0]�t!88�o�����|D�"���ɓ'���gǎ�yھ}{:D��ݫ�M�.]�l6SXX�޽{/���r�-�|>���HLL�j�����O?�Dtt4ݻw'((�3gΰu�V#�6�Lt�ܙ��x)--%55��6�DW��EDD�������#,,̘־}{ JKK�
Pxx86���g�r��	�N'$''T4��С6���Ktt4�{��`۽z����������Ǚ3gc��t����CBB�ׯ��˥�'5r��Q�����ݪU+<�E+�6��#G���w���7ߐ������			��6bbbe���lڴ������ILL䧟~���'  �>}��t�ԉΝ;��~���kRRR�֭;vl��BwDDD�Q���ݾ}{���'44Ԙ^yerǎ8�N�V+6���!C���'..����������~ *�"DEE�&11�h�w�^ z��I�N��ڵ+G���v�X,�o�Njj*&��h$R������Gjj*			U��s��<g�޽DFFҶm[�\���ɶmیu?~�:�|�r����C��ի��w<h�u+**"88��]�r��!%"""Rw������%22���8v��M�v퀊6�ǎ3捉��[�n_���� ��Oe%����!�M����v�J׮]�V��h֬Y���eee������r5IoBB999DFF�e����/�/00�N�:I@@ &�	��Jii�eן��_�t88�*�V�???l6V�������Ν;h4!R" """u"55���Hl6qqq����++?͚5�_�~�L&N�>Mjj*n���n�ɨ,���
QeBP��y333)**�`����1V���:v�=z��o߾F��%���r�k�.JJJ�x<�����3s)������ŕ:�������Թ����ݫW/�V+�ߝ��*W��������9}��1/T�(TYyiٲ�����Μ9c��v�ٳg��:p� W��*RS.����t�����K����',,�}�����CII	N���^��SZZ���@10    IDATr� 22����F;�������#^����4c��h����e̓������b�УG"""hӦM�����cǎO�v����SZZʡC�HJJ�]�v���Q\\l4/*--�2r�Hmٱc�w�������q:����Mvz��App0gϞ��}��|8p�.]�PRR��ӧ���"11�={�4�c�D@DD��IMM5:�BE3�s�&�y�f�w�NHHV��ЩS'�5kf̷s�N|>m۶%<<���\v��mt���{�n
���'44�f͚�p88y�$'N���:��x�x<���oܸ�޽{3r�H�n7uvN���`2��֭�������w��*C�66&I�l��;��%yP+�i�"""�MDD�O���2>���yAi:


�5��ng�T��7���{�# """"�)Q" """""JDDDDDD�������(%"""""�D@DDDDD�������Q" """""JDDDDDD�������(%"""""�D@DDDDD��������T"""���b��n�}����v���ظq#����<}���k׮DDD��/����^r}6���C�������d˖-�޽����"���X�c 2d:t ((���bv�������M����C}�>���/^ݢ>ڶ���\��""�(QZZZ��<v����Y�V���ذa�7o��r1l�0RRR(++�n����������r��Qcy��L�֭q8x�^��NBBBX�h���>�'NPXXp��W�J1\izC���r�c��n�JFFw�y'�O�&??�^�P��^nzC���~�Ng����"�t�W�S� �z�������S�NQZZ��ݻ),,�e˖�<�&55������?L���1��t�ԉM�6QZZJff&)))t��Ũ$]nz]�p��!���L
)++������r�7o^ob���6�����S" ""RO��ӧ�]�]�h������b�Z���5����p���+��7��O<����'�^/��71\�vB��Pߨ����H=d�X���{ٳggΜ��2>��'N WC++C�V�l6[��_�.6�!Űu�Vv��Ell,����~ԇ�u�!���}��tG@DD���s6�1b��u��]�:\.@����f3*:W�^�1T'��Cyy9EEE<x��J߾}�M����CC�>(�jU>��> V�\�����~~~<���`


p�\U�6DEE�[�4�.c����ń��֛�u�!���}P" """Wd2�>|8�Z�
�ٌ��&��J�����\�}�޽{���%%%��@LL����߿����*�+Mo1�l6���Chh(���t�ؑ.]����^ob���6�������T�K��^^�����X��""�(EDD��������tVa��BBB���\���u�عs' ���0���m۶�~�����l�u�]���_r���M�W��:1���V+#G��e˖X�V


ؽ{7?���E�w#b������������Z���v6n8Aŵ��?|��z��H��P5i�������(%"""""�D@DDDDD�������Q" """""JDDDDDD�������(%"""""�D@DDDDD��������)?���H�̝w�I߾}�ݻ7��ż���ܹS1� V��A�1x�`:w�L�-��|���r��!6l���p�\:��^0�H�UoV�y//ɃZQ\\�R�F)""�ӧO�h�χ��e˖u�Ov��1c�0j�(����LKOOg�����\C�4h�'O&::���eee1w�\~��G�FCAAA���T4�1���{�# ""�@��Ӈ��?�'QQQ�LB��e2�x�'x�ᇫ5ll,/��2�/f޼yx�^�K7��`ĈL�2������nݪ��?��O�N��������ܹsut.�0�,,""� ��g�y沕�u��)��(99����7W��o�[��sI�����\�s��<��ӘL�o3���CJJ�b�^(��'�x��3i�$�V��C>�n$5��������b�⼩����Mtc�!,,�|��Һuk�n7����n����Crr2����C�A�����T˨Q�����ּ������~��L�:����*����Z���Ht.���f���CU{~�ۭ� 	x����Zu��Iǡ	�P�����H=t��7^��Ͽb��MXXS�N��$ �Q�\j�1(�j�۷o�毫�5�|���V�

�7�`��:�8%"""R-=z�������WNQ1T�-��r]�׫W/fϞ͸q�tiJDDD�Z"##k4ppp�+K��Ҫ�)�6�L&���?p�M7�84������Y,���fذa����ȡ'ǎ����bP" """�b2���Y�СC���V� ++몖��_x��W7nw�}7w�u&L`�ܹ�:u�Z��ܹ��C#�����"""���������j/S\\̿���z3~zC�a���t�С��9s��^{�͛7_0---���4�,Y�o�[���?\��X.�Kǡ�ŠD@DDD�-##�������0u�T�?n<��[n�U�V���s��	6n�ȗ_~IQQ�b���?��_����9(##��������\q�.\HJJ
�g�������KII�qh�1�G/^ݢ>ڶ���\��""�(QZZZ��<�5?y6::�Z����x��'IKK��n���_�o߾�h�???�������O�>�5�#G�p�ĉ�R~9���2233����/�,���b�z�)N�<Y�}߾};����z�������o^u�$�K�#��Y��l6�E��"/%"""M2(..fĈW����f۶m�Sp/u����1d�RSS��Ȩ��k�1���q��q����f��<���o�o��m��V�}_�~=K�.eÆ���Ѯ];���������իux%0�H�f�x�y//ɃZQ\\��""�(EDDp���-���p:���@#������iӦ�%�9}�4�<�͚5c����N>���0a���u\�h�1 4oޜ|�ЦM���5���O>��}		�]�v�ٳGǡ�PPPP���v;7��b�%"""J��[o���_~���w���ڵkٹs'�������g���5Z��를���dɒ�vr��!�+y�ǘ0aB��w�K�7����i����%�ȦAP�4�O�>FRQVV��/�̼y�8x�q�'� <<�F�6�L���ï~�+,?��s��ac��J���?��}׹t}cP� ��F� �����w�%44��{�;vŤI����q������g�|ӧO�����!�s5�}׹t�b���F���N����&���K��|@RRV��ˎjS-Z�`͚5�^��!�s�����:��_厀�# ""R��߿� 0i�$BBB�d;��������]�R�;7���|����7�|�b����\%"""rQ��D[����_��#;wu/Y�D14��׹T?����y��QTTT����Oزe�bh�s�~�A����\B}5�|���|��wDFF��f��u9~���|�MV�Xq�ʵ!���_�R����#��g���h=G@DD���ix�sj�4�l61��n|�_O�(�����4P�~���l���=�4y11!8��$HDDDD��&&��_��S�:��N18��9�*9�ƚ�zk3f��[��x<�n�JLD�1�LX,,f��ɤB��χ�������x������[oMbڌ���; ���薭Gy덯	�?!�����c6����\^e���zq:�*3��%��'�ܴ{HN�xљwl?�+�\���R/ɃZ���j%((����*W�¹W����(--��r� ���$��3�|�U2�����+�X"зo;�|zC�v��L�:ʫ�\�ƍ�>T��f#,,�����M�ٌ�l�j�@���q:����U{,\�uy��0��������ȹ����c�����c�q�~���f����d2F�f̀��e���O���iժ �>}���L�m�Ɩ-[())������'::���"���t%M�F�P���j)�R" "rN�3�Ԛjw��g��5�X��9���{U4��j��l&22��� l6�F�� ((�˕����_�|��:}�sYY���x�^,��,00PM�j�����p�h���@1???&O�̭��ʱc�x������jp	�bP�%���@�*����'��k��jŮ�\�U"Pg�d"**��� Z�h�����رc��q��QfϞMnnn�����ԩS�3 r�]邀T_iii�H:t������ر#��� �ݻ�'�|��|?�0O<q��Ι3��˗0z�hF��+����w�M\\��RM;�s�=�I�&��W����(���>�SO~ʯ��+�����uV� <<�W_}��I @||<�g�&<<�����ߟ��00��m۶4��:ɉ���� t�֍5kְw�^.\H�.]�_�bh�1t�ԉ?�񏗜����.�n��Q���f�ѬY3l63f̸��|DDӧOgƌu�L�Y�f�i3$��m۶1b�JJJ�?>mڴ����w�fʔ)��~��	����_|��A�8q�D�7U/�����?������_�~���3�ɦF��s�N��?���ݻ�s�N}��������ܹ�T{��+���?			׼:t����8uW@��
dÆ<���t�ڕ6���Ns��h��Ν;�j�*���+�Ν���ë\�\�x1�\��1c��ꫯ*�p��S��?��N�<y�yC�R/��0��<��Ì9�֭[c�Z),,����_��O?�Ԙ��'���`��\�v�ݬ_�������X�~=������+����������_��׬Y���F
�j�j��Fd�ʕ���^v���x�6m�ġC�(**bӦM�8qBX�9JKK���&))��S��;�@aa!O<����Ui��T��<x0�-b���0��)%5���OW�|>���DFF��n��\Iyy9O=�����ﯔ��L�k:؏?�8&���},*; 0�V;ӿ֮][g�,00P��HT^^�ԩS���}/���͛��8u� ������DDD����GU�hTӎъ�i�о}{���?�w�^>���j-��T��w�����y�g(..&((�N�:o̷h�"���l��w�}�s�=��d����4�KOOgŊ,\��h�����^�zq���,Y���{Z�j�رc9x��E�q�ȑ�=����f3G���O?e����<���3�;v��+�]����}��z���۷����B��i$��~c�һ�ۨ���k�Z���o�Q�h׮&����V�^͒%K�����{�.]�p��A�,Y�ĉ	c�֭���d������'<<�}����+�4������*gee�c����b!""���+��C���Z�$%%��W_�*}��W,^���>�H1(����"""%11�}��QZZ�Ν;ٹs�1��Ç	#22���󑖖���>�#�<@nn.n���;��3�ЩS'fΜYe���������RTTt��{��?~< ;w����p��73k�,���kt��\����^ۮ�a�ZU4���s���{��c4�|ꩧx衇��+en����&O�Lbb"/��r�u�mۖ�3gRZZJ@@ ��vm۶�}�����H߾}�1c�'O�A�&L`Æ���W�o��&�8��ӊ�q�PYq>��\��ɰbP"pU>��^|�E:v��|���%--�-[��_��_F����oU�L�8���o~� 6n���O?����?��?>|8��s�~�))))�v����5k˖-�l6_th���h���{��ܹs�2e
�ƍ���3K�.����+�͛7��2�|
��111��׿`�֭L�:�����?�СC�뮻X�h�2�	䩧�������'))������o��g�1s�L��nz���f�hd5УG�M�@TT ����`3g��رc>�G}���


���6��-Z����UPM3��k�^��`ʔ)�9�:�bP"Pc+W����>�~�����H���i߾=��{/���o/ٳ�R׮]�/��ի���r�J�T�{n"p��i�-[�����Pݺu3���?��qgh߾=�WVς��ԩS'�p͚5�o��_�СC�ҥK�D ;;�;v p��1��� X�b G�*�f���+ 66��g6����f�0�|LBB�����瓞��_|��?��C�ch���� T<��w��w��j�2v�X�����΢E�j}�չW�f*�"���_0O~~�Um���`6�9{�l�?9��;�4ŬYDj��~D�͍\.�q����������m�6��+ηjժ*}<�b���7g��̙��\������w�f�֭dgg_pu���6�	

2n%�۷�χ�db���Y���˽��k̿w����޽{�z���fJJJx��i����z�dgg_ue�j�r��qZ�n]�eZ�oB���Ԇ���7vذa|��wx�^c�������DD��LϞ=�
������m�KKKY�n�1�ѣG���-�ԩS,Z��իW�h�"y����Y�jn����#?�YPuegg�p�B~���1r�H�u�Fzz:-[�$!!����*#�DYYlٲ�A��j�n޼�N����зG�	���f�ҥ<��C��ߟe˖�v������o���,HDD�T�o��m��F�n݈�� ((�3gΰk�.���*�֭[�ҥK2dQQQDEE�����;v�x���xL&�6��Zs����ѣ<��t�Ё֭[s��Y�l�������}uii)͛7租~�������Z)���b~��'%"R��z�-�?�ȑ#i׮f����Tc�PiXL&��٫�w��K�V����˗Ӻuk~���L�R�eZ�l��fc�ȑL�8�V����c�ʕU�Tզ��2u���j�QSV��Y"""j������t:iٲ�
\��*((��|v���N f�tޫ�wV-��������v�5 //������/�0��8p� _}�U�%��,""""��ZСC���éS�x������/��lyy9EEE�L&��fW+''�_|�N����"��-"""��iP�8&�����l������/ӹs��������o����Ά�s:��:uJ�(���4���i��\j$5�����Kyy9N��g�y���{����+.[\\�ܹsy��'�4	(++#''GI����7���"��^/999���a�������ꫯ��[HNN&..�����aaiiilܸ��7�r���}+**"//O��Dn`��.��5����������"�D@�����ٳӼysL&?�������bf��ٌ�j�j��YPVVF^^����`n��ͦ������T^^�D@D�H��y���`�Z	$00�͆�b���?^��ǃ����p�p8p�\:"��[��s��߸���VZZJ``���41���z��r�r�(,,Ta�4�*N�%W�8���M�Ʉ����p���HӐ���(""$(++��r��z�g��Uy���캗��b�d2QXXxݓ�q�Ng����;""H�B��L&���c��
		!((Ḧ́D)�χ��hp�8�������l܉(**��p����q�@Dv�����t:)--5$hH�m%"""��d2#U6�r��QTT�i��{��Ԡ�r]S"��T�m���"""�N*Ge��K���}�X,X,�ץl"P^�Q" ""r��pUi�����[^�{͉�ͦ6����{�m��0��m'��z�n���e`���i�Z�"	��\$����ۇ��#E�&q|����m  b ���V�����:1���W��  <Y� �H�T77������0�a�  IDAT��<>   h(I]]���NA��v��*'    B�r����E`�nB������k��s�(   P�b�з�7���A�x$/.~��n��l�R   *�f3�����^� %4�#��ӕB��E   (����L_>_��Gzנ��r�ѧ/5�/��   p MS-/���-���!�e����o��+}��?��nB   ��l6S����Ånn��o8U[�L�>�+^ҋ��z�V�^�Z���l6,}   <;I�h>���n�/��k��T����@� ��0 I�޽����"h��(�2�y���;k   �3��J�Di�j�����./���_`�A�\�^ x�z��߾ԛ7s-���DI£�  �td�k�δZmts���參�L+tu� �f�|�
�{���vmG{�V���gێW�ҏ�0K&��3�5�ڌV���$Z}��L�Ou� <��vU︑v��Eï��4���bl����m�@%Ŵu/�);3^5ioz��LL���d���37��X~m|���M߬�&���y+_IO�c� @Љ��ۇ��'��W����
�!�^�m*����.�Κ�*܊gP-B+A��Кϲ�Y�!��l��7��ѫf��Z`} +Y߭⛮_7�s/���x�8�U b߫��q�i��n8���H;���%e.e��dW�Z�v|X'y�P`��8��`:�6�vv��U��M�c��c ��U|�� �* ����ƕƛ�6- ;�Q���2��C ��6$�.�b�oR���T���,sײ��
X.yh[�U�G ��k��OuZ  b� "�sa ����5�����F+�Aw�3�
a�����=)��B�ph�R��� ��m��Zg�v" ���5��K����s�WMq{l\�b9�.X��Ż�8u=A��C�z|p�J��G�b�^g�4H��o ���I��
  ��tx\3 ��Nc�@ ���
�`p����t��t I$mY�>��A.yq������}�n@ 0^ 0�@p��)��,۵��-H�\a_�Z�q�A�"T���P݃��V�<~OM���-���5~�v�j�] x�  <�@�G�ֶ� ��w�

��>M�u��֟����]>T\�z ���?:� ����օ:�A x�����@�>� W�P�0�i����{��=��24���A�����ź�0 �D� <��uHd �~P@�P`��m(hT�W��B�EA�}ʰ�?G{;-�ï��� �9  ԭ�Z���'0IVh)(uV㶟���Zͧ�Vߓ0�S��5xOcT1Nk�:��� F�M @ @(�5?�}����j�ٷ����aT�I�~��4��t��|���4F ��   hX v�:$\S`�f����:���[�f.wk�����.g�{ �cI�    �b���b�`�����!�Ð݃&�؊u�=��_�|2�  �����p#���.D�b?��a���h8	�f��A�����9%���  ����(�s8e�    IEND�B`�