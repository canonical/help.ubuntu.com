<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" width="840" height="500" id="svg10075" version="1.1" ns1:version="0.92.4 5da689c313, 2019-01-14" ns2:docname="gs-datetime.svg">
  <ns0:defs id="defs10077">
    <ns0:linearGradient ns3:paint="gradient" id="RHEL7">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1;" offset="0" id="stop11074"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:1" offset="1" id="stop11076"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0;" offset="0" id="stop7012"/>
      <ns0:stop style="stop-color:#eeedec;stop-opacity:0" offset="1" id="stop7014"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#GNOME" id="linearGradient7064" gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" x1="-18.33782" y1="490.54935" x2="713.42853" y2="490.54935" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient5885" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720"/>
    </ns0:linearGradient>
    <ns0:linearGradient ns1:collect="always" ns4:href="#linearGradient5716" id="linearGradient17441" x1="29.089951" y1="11.772627" x2="33.971455" y2="9.7093649" gradientUnits="userSpaceOnUse"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop17445"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop17447"/>
    </ns0:linearGradient>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17453" ns4:href="#linearGradient5716" ns1:collect="always"/>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17455" ns4:href="#linearGradient5716" ns1:collect="always"/>
    <ns0:filter color-interpolation-filters="sRGB" ns1:collect="always" x="-0.10291173" width="1.2058235" y="-0.065432459" height="1.1308649" id="filter5601">
      <ns0:feGaussianBlur ns1:collect="always" stdDeviation="0.610872" id="feGaussianBlur5603"/>
    </ns0:filter>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17453-7" ns4:href="#linearGradient5716-4" ns1:collect="always" gradientTransform="matrix(1.0281734,0,0,1.0281734,637.14345,666.93836)"/>
    <ns0:linearGradient id="linearGradient5716-4">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop5718-1"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop5720-6"/>
    </ns0:linearGradient>
    <ns0:linearGradient y2="9.7093649" x2="33.971455" y1="11.772627" x1="29.089951" gradientUnits="userSpaceOnUse" id="linearGradient17455-1" ns4:href="#linearGradient5716-4" ns1:collect="always" gradientTransform="matrix(1.0281734,0,0,1.0281734,637.14345,666.93836)"/>
    <ns0:linearGradient id="linearGradient16929">
      <ns0:stop style="stop-color:#000000;stop-opacity:1;" offset="0" id="stop16931"/>
      <ns0:stop style="stop-color:#484848;stop-opacity:1;" offset="1" id="stop16933"/>
    </ns0:linearGradient>
  </ns0:defs>
  <ns2:namedview id="base" pagecolor="#eeeeec" bordercolor="#666666" borderopacity="1.0" ns1:pageopacity="1" ns1:pageshadow="2" ns1:zoom="1" ns1:cx="154.72357" ns1:cy="347.41188" ns1:document-units="px" ns1:current-layer="g4890" showgrid="false" borderlayer="true" ns1:showpageshadow="false" ns1:window-width="2560" ns1:window-height="1403" ns1:window-x="2560" ns1:window-y="0" ns1:window-maximized="1" width="0px" height="0px" fit-margin-top="0" fit-margin-left="0" fit-margin-right="0" fit-margin-bottom="0">
    <ns1:grid type="xygrid" id="grid17504" empspacing="5" visible="true" enabled="true" snapvisiblegridlinesonly="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g ns1:label="bg" ns1:groupmode="layer" id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true">
    <ns0:rect style="fill:url(#BLANK);" id="background" width="866" height="656" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g ns1:groupmode="layer" id="layer2" ns1:label="fg" transform="translate(0,-540)">
    <ns0:g id="g11020" transform="translate(-89,-139.36217)">
      <ns0:circle transform="translate(2,453.36217)" id="path11014" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;enable-background:accumulate" cx="120" cy="278" r="17"/>
      <ns0:text id="text11016" y="736.36218" x="122.29289" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="736.36218" x="122.29289" id="tspan11018" ns2:role="line" style="font-size:14px;line-height:1.25">3</ns0:tspan></ns0:text>
    </ns0:g>
    <ns0:g style="display:inline" id="g4890" transform="matrix(2.6833333,0,0,2.6833333,-1275.5101,-1072.8539)">
      <ns0:path style="display:inline;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-opacity:1" d="m 506.43234,611.75299 h 258.32299 c 2.21601,0 4,1.784 4,4 v 161.22982 h -4 -258.32299 -4 V 615.75299 c 0,-2.216 1.784,-4 4,-4 z" id="path5430" ns1:connector-curvature="0" ns2:nodetypes="sssccccss"/>
      <ns0:path ns1:connector-curvature="0" id="path5361" d="M 502.98343,630.36169 H 768.47408" style="display:inline;fill:none;stroke:#000000;stroke-width:1.01455009;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:nodetypes="cc"/>
      <ns0:path style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:xx-small;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#0c0000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1.3358984;marker:none;enable-background:new" id="path5375" d="m 756.48074,617.84776 h 0.74998 c 0.008,-9e-5 0.0156,-3.5e-4 0.0234,0 0.19121,0.008 0.38239,0.0964 0.51561,0.23437 l 1.71089,1.71088 1.73432,-1.71088 c 0.19921,-0.17287 0.335,-0.22912 0.51561,-0.23437 h 0.74998 v 0.74998 c 0,0.21484 -0.0258,0.41297 -0.1875,0.56248 l -1.71088,1.71089 1.68745,1.68745 c 0.14113,0.14112 0.21092,0.34008 0.21093,0.53905 v 0.74997 h -0.74998 c -0.19897,0 -0.39793,-0.0698 -0.53905,-0.21093 l -1.71088,-1.71089 -1.71089,1.71089 c -0.14112,0.14114 -0.34009,0.21093 -0.53905,0.21093 h -0.74998 v -0.74997 c 0,-0.19897 0.0698,-0.39793 0.21094,-0.53905 l 1.71088,-1.68745 -1.71088,-1.71089 c -0.15806,-0.14597 -0.22737,-0.35193 -0.21094,-0.56248 z" ns1:connector-curvature="0" ns2:nodetypes="ccccccccscccccscccscsccccc"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="669.13416" y="622.67847" id="text12012"><ns0:tspan ns2:role="line" id="tspan12014" x="669.13416" y="622.67847" style="font-size:5.21739101px;line-height:1.25">Datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:rect style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.7453416;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" id="rect9293" width="147.9503" height="93.540375" x="600.56281" y="634.97662" rx="0" ry="0"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="645.52429" id="text26176"><ns0:tspan ns2:role="line" id="tspan26178" x="610.1059" y="645.52429" style="font-size:5.21739101px;line-height:1.25">Automatisk datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:text id="text26182" y="652.2323" x="610.1059" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#babdb6;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="652.2323" x="610.1059" id="tspan26184" ns2:role="line" style="font-size:4.47205019px;line-height:1.25">Kräver internetåtkomst</ns0:tspan></ns0:text>
      <ns0:g id="g9286" transform="translate(-17.515526,-52.919256)">
        <ns0:g id="g3921" transform="matrix(0.37267081,0,0,0.37267081,493.07637,552.48134)" style="display:inline"/>
      </ns0:g>
      <ns0:rect width="5.9627328" height="5.9627328" x="-514.0741" y="617.82538" id="rect10837-5-8-1" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.3726708;marker:none;enable-background:new" transform="scale(-1,1)"/>
      <ns0:path d="m 512.58846,618.5707 h -0.37267 c -0.004,-4e-5 -0.008,-1.7e-4 -0.0117,0 -0.095,0.004 -0.19001,0.0479 -0.25621,0.11646 l -2.34696,2.13121 2.34698,2.13121 c 0.0701,0.0701 0.16899,0.10482 0.26786,0.10482 h 0.37267 v -0.37267 c 0,-0.0989 -0.0347,-0.19774 -0.10481,-0.26786 l -1.79962,-1.5955 1.79962,-1.59549 c 0.0785,-0.0725 0.11297,-0.17488 0.10481,-0.27951 z" ns1:connector-curvature="0" id="path10839-9-9-5" style="color:#bebebe;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:medium;line-height:normal;font-family:'Andale Mono';-inkscape-font-specification:'Andale Mono';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.66381985;marker:none;enable-background:new" ns2:nodetypes="ccsccccccccccc"/>
      <ns0:rect style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.3726708;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" id="rect15386" width="11.925466" height="11.925466" x="505.35666" y="615.02734" rx="1.4906832" ry="1.4906832"/>
      <ns0:path style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" d="M 600.56278,658.59462 H 748.51309" id="path9309" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
      <ns0:text id="text9311" y="667.88458" x="610.1059" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan y="667.88458" x="610.1059" id="tspan9313" ns2:role="line" style="font-size:5.21739101px;line-height:1.25">Automatisk tidszon</ns0:tspan></ns0:text>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#babdb6;fill-opacity:1;stroke:none" x="610.1059" y="674.59259" id="text9315"><ns0:tspan ns2:role="line" id="tspan9317" x="610.1059" y="674.59259" style="font-size:4.47205019px;line-height:1.25">Kräver internetåtkomst</ns0:tspan></ns0:text>
      <ns0:path ns1:connector-curvature="0" id="path9331" d="M 600.56278,680.95488 H 748.51309" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" ns2:nodetypes="cc"/>
      <ns0:rect ry="5.4602423" rx="5.4602423" y="665.09509" x="719.65601" height="10.92049" width="19.803892" id="rect939" style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:0.3726708"/>
      <ns0:circle r="4.4139271" cy="670.55194" cx="733.60791" id="circle941" style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:path ns2:nodetypes="cccccccc" id="path5567" d="M 97.089832,2.8483222 V 19.288556 l 3.712308,-3.623922 2.12132,4.331029 c 0.5196,1.171377 3.22086,0.229524 2.45278,-1.336875 l -2.09922,-4.496756 h 4.68458 z" style="color:#000000;display:block;overflow:visible;visibility:visible;opacity:0.6;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;filter:url(#filter5601);enable-background:accumulate" ns1:connector-curvature="0" transform="matrix(1.0281734,0,0,1.0281734,637.14345,666.93836)"/>
      <ns0:path style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17453-7);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1.02817345;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" d="m 736.42336,669.32166 v 16.90341 l 3.8169,-3.72602 2.18109,4.45305 c 0.53423,1.20438 3.3116,0.23599 2.52188,-1.37454 l -2.15837,-4.62345 h 4.81656 z" id="path5565" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
      <ns0:path ns2:nodetypes="cccccccc" id="path6242" d="m 736.42336,669.32166 v 16.90341 l 3.8169,-3.72602 2.18109,4.45305 c 0.53423,1.20438 3.3116,0.23599 2.52188,-1.37454 l -2.15837,-4.62345 h 4.81656 z" style="color:#000000;display:block;overflow:visible;visibility:visible;fill:url(#linearGradient17455-1);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1.02817345;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:accumulate" ns1:connector-curvature="0"/>
      <ns0:path style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" d="M 600.56278,703.31514 H 748.51309" id="path9337" ns1:connector-curvature="0" ns2:nodetypes="cc"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="694.71686" id="text9333"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" ns2:role="line" id="tspan9335" x="610.1059" y="694.71686">Datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:text id="text9341" y="694.71686" x="740.54083" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" y="694.71686" x="740.54083" id="tspan9343" ns2:role="line">1 september 2015, 09:51</ns0:tspan></ns0:text>
      <ns0:text id="text9345" y="717.82251" x="610.1059" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" y="717.82251" x="610.1059" id="tspan9347" ns2:role="line">Tidszon</ns0:tspan></ns0:text>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="740.54083" y="717.82251" id="text9349"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" ns2:role="line" id="tspan9351" x="740.54083" y="717.82251">CEST (Stockholm, Sverige)</ns0:tspan></ns0:text>
      <ns0:rect ry="0" rx="0" y="742.30591" x="600.56281" height="23.478262" width="147.9503" id="rect9353" style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.7453416;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate"/>
      <ns0:text xml:space="preserve" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:start;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:start;display:inline;fill:#000000;fill-opacity:1;stroke:none" x="610.1059" y="756.2077" id="text9355"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" ns2:role="line" id="tspan9357" x="610.1059" y="756.2077">Tidsformat</ns0:tspan></ns0:text>
      <ns0:rect style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:0.37267077;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" id="rect9363" width="38.341366" height="12.298138" x="702.89008" y="747.73126" rx="1.0248625" ry="1.0248625"/>
      <ns0:text id="text9359" y="755.83502" x="727.87006" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell, Normal';text-align:end;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:end;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" y="755.83502" x="727.87006" id="tspan9361" ns2:role="line">24-timmars</ns0:tspan></ns0:text>
      <ns0:path style="color:#000000;clip-rule:nonzero;display:inline;overflow:visible;visibility:visible;opacity:1;isolation:auto;mix-blend-mode:normal;color-interpolation:sRGB;color-interpolation-filters:linearRGB;solid-color:#000000;solid-opacity:1;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0.3726708;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal;color-rendering:auto;image-rendering:auto;shape-rendering:auto;text-rendering:auto;enable-background:accumulate" d="m 737.50428,752.6939 -1.96993,1.96993 -1.96993,-1.96993 z" id="rect9365" ns1:connector-curvature="0" ns2:nodetypes="cccc"/>
      <ns0:text id="text946" y="622.67847" x="541.68079" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#000000;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan style="font-size:5.21739101px;line-height:1.25" y="622.67847" x="541.68079" id="tspan944" ns2:role="line">Detaljer</ns0:tspan></ns0:text>
      <ns0:rect transform="scale(-1,1)" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:0.3726708;marker:none;enable-background:new" id="rect948" y="617.82538" x="-575.56482" height="5.9627328" width="5.9627328"/>
      <ns0:rect ry="1.4906832" rx="1.4906832" y="615.02734" x="566.84741" height="11.925466" width="11.925466" id="rect952" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:0.3726708;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate"/>
      <ns0:g ns1:label="open-menu" id="g7352" transform="matrix(0.37267081,0,0,0.37267081,562.5214,515.34088)" style="display:inline;enable-background:new">
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" id="rect7354" width="16" height="16" x="20" y="276"/>
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7356" width="9.9996014" height="2.0002136" x="23.000198" y="278.99979"/>
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7358" width="9.9996014" height="2.0002136" x="23.000198" y="282.99979"/>
        <ns0:rect style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#2e3436;fill-opacity:1;stroke:none;stroke-width:1;marker:none" id="rect7360" width="9.9996014" height="2.0002136" x="23.000198" y="286.99979"/>
      </ns0:g>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#000000;fill-opacity:1;stroke:none;stroke-width:5.96273279;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7822" width="79.006218" height="17.142857" x="502.923" y="646.15674"/>
      <ns0:g ns1:label="preferences-system-time" id="g24827" transform="matrix(0.37267081,0,0,0.37267081,440.68702,454.60394)" style="fill:#ffffff;enable-background:new">
        <ns0:circle style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#ffffff;stroke-width:2.15384626;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" id="path24839" transform="matrix(0.92857143,0,0,0.92857143,198.85734,238.42857)" cx="-9" cy="321" r="7"/>
        <ns0:path style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#f7f7f7;stroke-width:1;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;enable-background:new" d="m -13.5625,316.46875 3.111031,3.04475 m 0.0029,-0.0135 h 2.948604" id="path25609" ns1:original-d="m -13.5625,316.46875 3.111031,3.04475 m 0.0029,-0.0135 h 2.948604" ns1:connector-curvature="0" transform="translate(201.0002,217)" ns2:nodetypes="cccc"/>
      </ns0:g>
      <ns0:text id="text7826" y="656.21881" x="536.0907" style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;display:inline;fill:#ffffff;fill-opacity:1;stroke:none" xml:space="preserve"><ns0:tspan style="font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;font-size:5.21739101px;line-height:1.25;font-family:Cantarell;-inkscape-font-specification:Cantarell;fill:#ffffff" y="656.21881" x="536.0907" id="tspan7824" ns2:role="line">Datum &amp; tid</ns0:tspan></ns0:text>
      <ns0:path style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:#000000;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" d="m 582.12691,611.30064 v 164.9182" id="path7828" ns1:connector-curvature="0"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7830" width="17.888199" height="3.3540373" x="521.92926" y="636.83997"/>
      <ns0:rect y="670.38031" x="521.92926" height="3.3540373" width="17.888199" id="rect7832" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:rect style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="rect7834" width="17.888199" height="3.3540373" x="521.92926" y="685.28717"/>
      <ns0:rect y="685.28717" x="544.28955" height="3.3540373" width="28.695652" id="rect7836" style="opacity:1;vector-effect:none;fill:#070707;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="path7840" cx="511.711" cy="638.71655" r="4.2555118"/>
      <ns0:circle r="4.2555118" cy="672.62958" cx="511.711" id="circle7842" style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal"/>
      <ns0:circle style="opacity:1;vector-effect:none;fill:#c0bfbc;fill-opacity:1;stroke:none;stroke-width:0.3726708;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="circle7844" cx="511.711" cy="686.79108" r="4.2555118"/>
    </ns0:g>
    <ns0:rect style="display:inline;fill:#000000;fill-opacity:1;stroke:none;stroke-width:1" id="rect3923" width="53.140442" height="29.303314" x="655.56671" y="645.81787" rx="14.65165" ry="14.65165"/>
    <ns0:circle style="opacity:1;vector-effect:none;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:16;stroke-linecap:round;stroke-linejoin:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-dashoffset:0;stroke-opacity:1;marker:none;marker-start:none;marker-mid:none;marker-end:none;paint-order:normal" id="path915" cx="693.00433" cy="660.46039" r="11.844038"/>
  </ns0:g>
</ns0:svg>
