<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Nätverkstermer &amp; -tips</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Nätverkstermer &amp; -tips</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="net-proxy.html" title="Definiera proxyinställningar"><span class="title">Definiera proxyinställningar</span><span class="linkdiv-dash"> — </span><span class="desc">En proxy filtrerar webbsidor som du tittar på, oftast av kontroll- eller säkerhetssyfte.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-findip.html" title="Hitta din IP-adress"><span class="title">Hitta din IP-adress</span><span class="linkdiv-dash"> — </span><span class="desc">Att känna till din IP-adress kan hjälpa dig upptäcka nätverksproblem.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-security-tips.html" title="Trygghet på internet"><span class="title">Trygghet på internet</span><span class="linkdiv-dash"> — </span><span class="desc">Allmänna tips när du använder internet</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="net-what-is-ip-address.html" title="Vad är en IP-adress?"><span class="title">Vad är en IP-adress?</span><span class="linkdiv-dash"> — </span><span class="desc">En IP-adress är som ett telefonnummer för din dator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="net-macaddress.html" title="Vad är en MAC-adress?"><span class="title">Vad är en MAC-adress?</span><span class="linkdiv-dash"> — </span><span class="desc">Den unika identifieraren som tilldelats din nätverkshårdvara.</span></a></div>
</div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a><span class="desc"> — <span class="link"><a href="net-wireless.html" title="Trådlös anslutning">Trådlöst</a></span>, <span class="link"><a href="net-wired.html" title="Trådbunden anslutning">trådbundet</a></span>, <span class="link"><a href="net-problem.html" title="Nätverksproblem">anslutnings-problem</a></span>, <span class="link"><a href="net-browser.html" title="Webbläsare">webbnavigering</a></span>, <span class="link"><a href="net-email.html" title="E-post &amp; e-postmjukvara">e-postkonton</a></span>, <span class="link"><a href="net-chat.html" title="Chatt &amp; sociala medier">snabbmeddelanden</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless.html" title="Trådlös anslutning">Trådlös anslutning</a><span class="desc"> — <span class="link"><a href="net-wireless-connect.html" title="Anslut till ett trådlöst nätverk">Anslut till trådlöst nätverk</a></span>, <span class="link"><a href="net-wireless-hidden.html" title="Anslut till ett dolt, trådlöst nätverk">Dolda nätverk</a></span>, <span class="link"><a href="net-wireless-edit-connection.html" title="Redigera en trådlös anslutning">Redigera anslutningsinställningar</a></span>, <span class="link"><a href="net-wireless-disconnecting.html" title="Varför kopplar mitt trådlösa nätverk ner hela tiden?">Nedkoppling</a></span>...</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
