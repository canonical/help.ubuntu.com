<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Bläddra bland filer och mappar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Bläddra bland filer och mappar</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Använd filhanteraren <span class="app">Filer</span> för att bläddra bland och organisera filerna på din dator. Du kan också använda programmet till att hantera filer på lagringsenheter (t.ex. externa hårddiskar), på <span class="link"><a href="nautilus-connect.html" title="Bläddra bland filer på en server eller nätverksdelning">filservrar</a></span>, och i delade mappar på ett nätverk.</p>
<p class="p">För att starta filhanteraren, öppna <span class="app">Filer</span> i <span class="gui">programstartaren</span>. Du kan också söka efter filer och mappar med <span class="gui">Dash</span> på samma sätt som du <span class="link"><a href="unity-dash-intro.html#dash-home" title="Search everything from the Dash home">söker efter program</a></span>. De visas sedan under rubriken <span class="gui">Filer och mappar</span>.</p>
</div>
<div id="files-view-folder-contents" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Utforska mappars innehåll</span></h2></div>
<div class="region"><div class="contents">
<p class="p">I filhanteraren, dubbelklicka på en mapp för att visa dess innehåll, och dubbelklicka på en fil för att öppna den med det förvalda programmet för den filen. Du kan också högerklicka på en mapp och öppna den i en ny flik eller ett nytt fönster.</p>
<p class="p"><span class="em">Sökvägsraden</span> ovanför listan över filer och mappar visar dig vilken mapp du tittar på, inklusive överstående mappar för den aktuella mappen. Klicka på en överstående mapp i sökvägsraden för att gå till den mappen. Högerklicka på en av mapparna i raden för att öppna den i en ny flik eller nytt fönster, kopiera eller flytta den, eller kom åt dess egenskaper.</p>
<p class="p">Om du snabbt vill gå till en fil i mappen du visar, börja skriva in filens namn. En sökruta kommer visas överst i fönstret, och den första filen som matchar din sökning kommer markeras. Tryck på neråtpilen eller rulla med mushjulet för att gå till nästa fil som matchar din sökning.</p>
<p class="p">Du kan snabbt komma åt vanliga platser från <span class="em">sidoraden</span>. Om du inte ser sidoraden, klicka på <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="nerknappen"></span></span> i verktygsraden och välj <span class="gui">Visa sidoraden</span>. Du kan lägga till bokmärken till mappar som du använder ofta, så visas de i sidoraden. Använd menyn <span class="gui">Bokmärken</span> för att göra det, eller dra en mapp till sidoraden.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files-copy.html" title="Kopiera eller flytta filer och mappar">Kopiera eller flytta filer och mappar</a><span class="desc"> — Kopiera eller flytta objekt till en ny mapp.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
