<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Use different speakers or headphones</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="media.html#sound" title="Grundinställningar ljud">Ljud</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Use different speakers or headphones</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">You can use external speakers or headphones with your computer. Speakers
  usually either connect using a circular TRS (<span class="em">tip, ring, sleeve</span>) plug
  or with USB.</p>
<p class="p">If your speakers or headphones have a TRS plug, plug it into the appropriate
  socket on your computer. Most computers have two sockets: one for microphones
  and one for speakers. Look for a picture of headphones next to the socket.
  Speakers or headphones plugged into a TRS socket will usually be used by default.
  If not, see the instructions below for selecting the default device.</p>
<p class="p">Some computers support multi-channel output for surround sound. This usually
  uses multiple TRS jacks, which are often color-coded. If you are unsure which
  plugs go in which sockets, you can test the sound output in the sound settings.
  Click the <span class="gui">sound menu</span> on the <span class="gui">menu bar</span> then click
  <span class="gui">Sound Settings</span>. Select your speakers in the list
  of devices, then click <span class="gui">Test Sound</span>. In the pop-up window, click the
  button for each speaker. Each button will speak its position only to the channel
  corresponding to that speaker.</p>
<p class="p">If you have USB speakers or headphones, or analog headphones plugged
  into a USB sound card, plug them into any USB port. USB speakers act as
  separate audio devices, and you may have to specify which speakers to
  use by default.</p>
<div class="steps"><div class="inner">
<div class="title title-steps"><h2><span class="title">Select a default audio input device</span></h2></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Click the <span class="gui">sound menu</span> on the <span class="gui">menu bar</span> and select <span class="gui">Sound Settings</span>.</p></li>
<li class="steps"><p class="p">On the <span class="gui">Output</span> tab, select the device in the list of devices.</p></li>
</ol></div>
</div></div>
<p class="p">If you don't see your device on the <span class="gui">Output</span> tab, check the
  <span class="gui">Hardware</span> tab. Select your device and try different profiles.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="media.html#sound" title="Grundinställningar ljud">Grundinställningar ljud</a><span class="desc"> — <span class="link"><a href="sound-volume.html" title="Change the sound volume">Volym</a></span>, <span class="link"><a href="sound-usespeakers.html" title="Use different speakers or headphones">högtalare och hörlurar</a></span>, <span class="link"><a href="sound-usemic.html" title="Använd en annan mikrofon">mikrofoner</a></span>...</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="sound-usemic.html" title="Använd en annan mikrofon">Använd en annan mikrofon</a><span class="desc"> — Use an analog or USB microphone and select a default input device.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
