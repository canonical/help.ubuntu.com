<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vad betyder ikonerna i systemraden?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 25.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html.sv" title="Ditt skrivbord">Skrivbord</a> › <a class="trail" href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Vad betyder ikonerna i systemraden?</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Denna sida förklarar innebörden av ikonerna som finns i det övre högra hörnet av skärmen. Mer specifikt förklaras de olika varianterna av ikoner som erbjuds av systemet.</p>
<div role="navigation" class="links sectionlinks"><div class="inner"><div class="region"><ul>
<li class="links "><a href="status-icons.html.sv#universalicons" title="Hjälpmedelsikoner">Hjälpmedelsikoner</a></li>
<li class="links "><a href="status-icons.html.sv#audioicons" title="Ljudikoner">Ljudikoner</a></li>
<li class="links "><a href="status-icons.html.sv#batteryicons" title="Batteriikoner">Batteriikoner</a></li>
<li class="links "><a href="status-icons.html.sv#bluetoothicons" title="Bluetooth-ikoner">Bluetooth-ikoner</a></li>
<li class="links "><a href="status-icons.html.sv#networkicons" title="Nätverksikoner">Nätverksikoner</a></li>
<li class="links "><a href="status-icons.html.sv#othericons" title="Övriga ikoner">Övriga ikoner</a></li>
</ul></div></div></div>
</div>
<section id="universalicons"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Hjälpmedelsikoner</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-accessibility.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Låter dig snabbt växla diverse hjälpmedelsinställningar.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-pointer.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar klicktypen som kommer att ske vid användning av uppehållsklick.</p></td>
</tr>
</table></div></div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="a11y.html.sv" title="Hjälpmedel">Lär dig mer om hjälpmedel.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="a11y-dwellclick.html.sv" title="Simulera klick genom att sväva ovanför">Lär dig mer om uppehållsklick.</a></span></p></li>
</ul></div></div></div>
</div></div>
</div></section><section id="audioicons"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Ljudikoner</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-audio-volume.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar volymen för högtalarna eller hörlurarna.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-audio-volume-muted.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Högtalarna eller hörlurarna är tystade.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-microphone-sensitivity.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar mikrofonens känslighet.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-microphone-sensitivity-muted.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Mikrofonen är tystad.</p></td>
</tr>
</table></div></div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="sound-volume.html.sv" title="Ändra ljudvolymen">Lär dig mer om ljudvolym.</a></span></p></li></ul></div></div></div>
</div></div>
</div></section><section id="batteryicons"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Batteriikoner</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-battery-charging.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar batterinivån då batteriet laddas.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-battery-level-100-charged.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är fulladdat och laddas.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-battery-discharging.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar batterinivån då batteriet inte laddas.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-battery-level-100.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Batteriet är fulladdat och laddas inte.</p></td>
</tr>
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-system-shutdown.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Strömikon som visas på system utan något batteri.</p></td>
</tr>
</table></div></div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="power-status.html.sv" title="Kontrollera batteristatus">Lär dig mer om batteristatus.</a></span></p></li></ul></div></div></div>
</div></div>
</div></section><section id="bluetoothicons"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Bluetooth-ikoner</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-airplane-mode.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Flygplansläge är på. Bluetooth är inaktiverat när flygplansläge är på.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-bluetooth-active.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">En Bluetooth-enhet har parats ihop och används. Denna ikon visas endast när det finns en aktiv enhet, inte bara för att Bluetooth är aktiverat.</p></td>
</tr>
</table></div></div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="net-wireless-airplane.html.sv" title="Stäng av trådlöst (flygplansläge)">Lär dig mer om flygplansläge.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="bluetooth.html.sv" title="Bluetooth">Lär dig mer om Bluetooth.</a></span></p></li>
</ul></div></div></div>
</div></div>
</div></section><section id="networkicons"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Nätverksikoner</span></h2></div>
<div class="region">
<div class="contents pagewide">
<div class="table"><div class="inner">
<div class="title title-table"><h3><span class="title">Trådlösa anslutningar (Wi-Fi)</span></h3></div>
<div class="region"><table class="table">
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-airplane-mode.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Flygplansläge är på. Trådlöst nätverk är avslaget när flygplansläge är på.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-network-wireless-acquiring.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluter till ett trådlöst nätverk.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-wireless-signal.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar styrkan hos en trådlös nätverksanslutning.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-network-wireless-signal-none.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådlöst nätverk, men det finns ingen signal.</p></td>
</tr>
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-network-wireless-connected.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådlöst nätverk. Denna ikon visas endast om signalstyrkan inte kan avgöras, såsom vid anslutning till ad hoc-nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-network-wireless-no-route.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådlöst nätverk, men det finns ingen väg till internet. Detta kan bero på en felkonfiguration av ditt nätverk, eller så kan det vara beroende på ett problem hos din internetleverantör.</p></td>
</tr>
</table></div>
</div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="net-wireless-airplane.html.sv" title="Stäng av trådlöst (flygplansläge)">Lär dig mer om flygplansläge.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="net-wireless-connect.html.sv" title="Anslut till ett trådlöst nätverk">Lär dig mer om trådlösa nätverk.</a></span></p></li>
</ul></div></div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h3><span class="title">Mobilnätverk (mobilt bredband)</span></h3></div>
<div class="region"><table class="table">
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-airplane-mode.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Flygplansläge är på. Mobilnätverk är avslaget när flygplansläge är på.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-network-cellular-acquiring.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluter till ett mobilnätverk.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-cellular-signal.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar styrkan hos en mobilnätverksanslutning.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-network-cellular-signal-none.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett mobilnätverk, men det finns ingen signal.</p></td>
</tr>
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-network-cellular-connected.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett mobilnätverk. Denna ikon visas endast om signalstyrkan inte kan avgöras, såsom vid anslutning över Bluetooth. Om signalstyrkan kan avgöras visas i stället en signalstyrkeikon.</p></td>
</tr>
</table></div>
</div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="net-wireless-airplane.html.sv" title="Stäng av trådlöst (flygplansläge)">Lär dig mer om flygplansläge.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="net-mobile.html.sv" title="Anslut till mobilt bredband">Lär dig mer om mobilnätverk.</a></span></p></li>
</ul></div></div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h3><span class="title">Trådbundna anslutningar</span></h3></div>
<div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-wired-acquiring.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluter till ett trådbundet nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-wired.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådbundet nätverk.</p></td>
</tr>
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-wired-disconnected.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ej ansluten till nätverket.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-wired-no-route.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett trådbundet nätverk, men det finns ingen väg till internet. Detta kan bero på en felkonfiguration av ditt nätverk, eller så kan det vara beroende på ett problem hos din internetleverantör.</p></td>
</tr>
</table></div>
</div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="net-wired-connect.html.sv" title="Anslut till ett trådbundet nätverk (Ethernet)">Lär dig mer om trådbundna nätverk.</a></span></p></li></ul></div></div></div>
<div class="table"><div class="inner">
<div class="title title-table"><h3><span class="title">VPN (virtuellt privat nätverk)</span></h3></div>
<div class="region"><table class="table">
<tr>
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-vpn-acquiring.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluter till ett virtuellt privat nätverk.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image"><div class="inner"><img src="figures/topbar-network-vpn.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluten till ett virtuellt privat nätverk.</p></td>
</tr>
</table></div>
</div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact"><li class="list"><p class="p"><span class="link"><a href="net-vpn-connect.html.sv" title="Anslut till ett VPN">Lär dig mer om virtuella privata nätverk.</a></span></p></li></ul></div></div></div>
</div>
<section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links seealsolinks"><div class="inner">
<div class="title"><h3><span class="title">Se även</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlösa nätverk</a><span class="desc"> — Anslut till trådlösa nätverk, inklusive dolda nätverk och nätverk består av en surfzon från en telefon.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
</div></section><section id="othericons"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Övriga ikoner</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="table"><div class="inner"><div class="region"><table class="table">
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-input-method.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Indikerar tangentbordslayouten eller inmatningsmetoden som för närvarande används. Klicka för att välja en annan layout. Menyn för tangentbordslayout visas endast om du har flera inmatningsmetoder konfigurerade.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-find-location.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ett program har för närvarande åtkomst till din plats. Du kan inaktivera platsåtkomst från menyn.</p></td>
</tr>
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-night-light.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Nattbelysning har ändrat färgtemperaturen för skärmen för att reducera trötthet i ögonen. Du kan tillfälligt inaktivera nattbelysning från menyn.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-media-record.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Du spelar för närvarande in en inspelning av hela skärmen.</p></td>
</tr>
<tr>
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-screen-shared.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ett program delar för närvarande skärmen eller ett annat fönster.</p></td>
</tr>
<tr class="shade">
<td><div class="media media-image floatend"><div class="inner"><img src="figures/topbar-thunderbolt-acquiring.svg" class="media media-block" alt=""></div></div></td>
<td><p class="p">Ansluter till en Thunderbolt-enhet, såsom en docka.</p></td>
</tr>
</table></div></div></div>
<div class="list"><div class="inner"><div class="region"><ul class="list compact">
<li class="list"><p class="p"><span class="link"><a href="keyboard-layouts.html.sv" title="Använd alternativa tangentbordslayouter">Lär dig mer om tangentbordslayouter.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="privacy-location.html.sv" title="Kontrollera platstjänster">Lär dig mer om sekretess och platstjänster.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="display-night-light.html.sv" title="Justera färgtemperaturen för din skärm">Lär dig mer om nattbelysning och färgtemperatur.</a></span></p></li>
<li class="list"><p class="p"><span class="link"><a href="screen-shot-record.html.sv" title="Skärmbilder och skärminspelningar">Lär dig mer om skärmbilder och skärminspelningar.</a></span></p></li>
</ul></div></div></div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html.sv#apps" title="Program och fönster">Program och fönster</a></li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
