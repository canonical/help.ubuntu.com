<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Fotolinsen</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="unity-dash-intro.html" title="Hitta program, filer, musik med mera med Snabbstartspanelen">Hitta program, filer, musik med mera med Snabbstartspanelen</a> › <a class="trail" href="unity-dash-intro.html#dash-lenses" title="Vyer">Vyer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Fotolinsen</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Fotolinsen är den femte linsen efter Snabbstartspanelens hem i <span class="gui">linsraden</span> och visas som en kamera. Fotolinsern låter dig komma åt foton på din dator eller från <span class="link"><a href="accounts.html" title="Nätkonton">Online-konton</a></span> som Facebook eller Google Picasa.</p>
<p class="p">Du kan använda <span class="keyseq"><span class="key"><kbd>Super</kbd></span>+<span class="key"><kbd>C</kbd></span></span> för att öppna Snabbstartspanelen direkt på fotolinsen.</p>
</div>
<div id="dash-apps-previews" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Förhandsvisningar</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Högerklicka på ett sökresultat för att öppna en <span class="gui">förhandsgranskning</span> med mer information om bilden och en större miniatyrbild.</p>
<p class="p">För foton som finns lagrade på din dator kan du välja att öppna, skriva ut, visa, eller skicka dem via e-post.</p>
</div></div>
</div></div>
<div id="dash-apps-filters" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Filter</span></h2></div>
<div class="region"><div class="contents"><p class="p">Klicka på <span class="gui">Filtrera resultat</span> för att filtrera efter vilket datum bilden togs, eller efter källa.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="unity-dash-intro.html#dash-lenses" title="Vyer">Vyer</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links "><a href="unity-dash-intro.html#dash-lenses" title="Vyer">Vyer</a></li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
