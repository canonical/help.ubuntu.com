<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>På/av &amp; batteri</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">På/av &amp; batteri</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="power-batterylife.html" title="Använd mindre ström och förbättra batteridriftstiden"><span class="title">Använd mindre ström och förbättra batteridriftstiden</span><span class="linkdiv-dash"> — </span><span class="desc">Tips på hur du reducerar din dators strömförbrukning.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-batteryoptimal.html" title="Få ut det mesta ur din bärbara dators batteri"><span class="title">Få ut det mesta ur din bärbara dators batteri</span><span class="linkdiv-dash"> — </span><span class="desc">Tips så som “Låt inte batteriet bli för lågt“</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-hibernate.html" title="Hur försätter jag min dator i viloläge?"><span class="title">Hur försätter jag min dator i viloläge?</span><span class="linkdiv-dash"> — </span><span class="desc">Viloläge är inaktiverat som standard eftersom det saknar bra stöd.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-exit.html" title="Logga ut, stäng av, växla användare"><span class="title">Logga ut, stäng av, växla användare</span><span class="linkdiv-dash"> — </span><span class="desc">Lär dig hur du lämnar ditt användarkonto, genom att logga ut, byta användare, och så vidare.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-suspend.html" title="Vad händer när jag försätter min dator i vänteläge?"><span class="title">Vad händer när jag försätter min dator i vänteläge?</span><span class="linkdiv-dash"> — </span><span class="desc">Vänteläge försätter din dator i ett strömsparläge där den drar mindre ström.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-closelid.html" title="Varför stängs min dator av när jag stänger locket?"><span class="title">Varför stängs min dator av när jag stänger locket?</span><span class="linkdiv-dash"> — </span><span class="desc">Bärbara datorer försätts i strömsparläge när du stänger locket för att spara ström.</span></a></div>
</div></div></div></div>
<div id="battery" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Batteriinställningar</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="power-batteryestimate.html" title="Den uppskattade batteridriftstiden är fel"><span class="title">Den uppskattade batteridriftstiden är fel</span><span class="linkdiv-dash"> — </span><span class="desc">Batteridriftstiden som visas när du klickar på <span class="gui">batteriikonen</span> är en uppskattning.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-batterywindows.html" title="Varför har jag mindre batteridriftstid än jag hade i Windows/Mac OS?"><span class="title">Varför har jag mindre batteridriftstid än jag hade i Windows/Mac OS?</span><span class="linkdiv-dash"> — </span><span class="desc">Justeringar från tillverkaren och olika batteridriftsuppskattningar kan vara orsaken till detta problem.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-lowpower.html" title="Varför stängde min dator av/försattes i vänteläge när batteriet gick ner till 10%?"><span class="title">Varför stängde min dator av/försattes i vänteläge när batteriet gick ner till 10%?</span><span class="linkdiv-dash"> — </span><span class="desc">Att låta batteriet laddas ur helt är dåligt för batteriet.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="power-whydim.html" title="Varför tonas min skärm ner efter ett tag?"><span class="title">Varför tonas min skärm ner efter ett tag?</span><span class="linkdiv-dash"> — </span><span class="desc">När din bärbara dator körs på batteriström kommer skärmen bli mörkare när datorn inte används för att spara ström.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="power-batteryslow.html" title="Varför är min bärbara dator så långsam när den kör på batteri?"><span class="title">Varför är min bärbara dator så långsam när den kör på batteri?</span><span class="linkdiv-dash"> — </span><span class="desc">Vissa bärbara datorer kör avsiktligt saktare när de kör på batteri.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="problems" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Problem</span></h2></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region"><ul>
<li class="links "><a href="power-constantfan.html" title="Den bärbara datorns fläkt kör alltid">Den bärbara datorns fläkt kör alltid</a></li>
<li class="links "><a href="power-batterybroken.html" title="Ett felmeddelande visar att mitt batteri har låg kapacitet">Ett felmeddelande visar att mitt batteri har låg kapacitet</a></li>
<li class="links "><a href="power-nowireless.html" title="Jag har inget trådlöst nätverk när jag väcker datorn">Jag har inget trådlöst nätverk när jag väcker datorn</a></li>
<li class="links "><a href="power-othercountry.html" title="Kommer min dator att fungera med ett strömaggregat i ett annat land?">Kommer min dator att fungera med ett strömaggregat i ett annat land?</a></li>
<li class="links "><a href="power-hotcomputer.html" title="Min dator blir väldigt varm">Min dator blir väldigt varm</a></li>
<li class="links "><a href="power-willnotturnon.html" title="Min dator vill inte starta">Min dator vill inte starta</a></li>
<li class="links "><a href="display-dimscreen.html" title="Ställ in skärmens ljusstyrka">Ställ in skärmens ljusstyrka</a></li>
<li class="links "><a href="power-suspendfail.html" title="Varför återstartar inte min dator efter att jag har försatt den i vänteläge?">Varför återstartar inte min dator efter att jag har försatt den i vänteläge?</a></li>
</ul></div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h3><span class="title">Mer information</span></h3></div>
<div class="region"><ul><li class="links "><a href="hardware.html#problems" title="Vanliga problem">Hårdvaruproblem</a></li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="prefs.html" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html" title="Användarkonton">användarkonton</a></span>…</span>
</li>
<li class="links ">
<a href="hardware.html" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a><span class="desc"> — <span class="link"><a href="hardware.html#problems" title="Vanliga problem">Hårdvaruproblem</a></span>, <span class="link"><a href="printing.html" title="Utskrifter">skrivare</a></span>, <span class="link"><a href="power.html" title="På/av &amp; batteri">på/av-funktioner</a></span>, <span class="link"><a href="color.html" title="Hantera färginställningar">färginställningar</a></span>, <span class="link"><a href="bluetooth.html" title="Bluetooth">Bluetooth</a></span>, <span class="link"><a href="disk.html" title="Hårddiskar &amp; lagring">hårddiskar</a></span>…</span>
</li>
</ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
