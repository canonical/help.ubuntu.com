<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Snabbmeddelanden på Ubuntu</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-chat.html" title="Chatt &amp; sociala medier">Chatt &amp; sociala medier</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Snabbmeddelanden på Ubuntu</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Med programmet <span class="app">Empathy</span> kan du chatta med folk på nätet och med vänner och kollegor som använder Google Talk, AIM, Windows Live, och många andra chattprogram. Med en mikrofon eller webbkamera kan du också föra ljud- eller videosamtal.</p>
<p class="p">Empathy är inte installerat i Ubuntu som standard, men du kan <span class="link"><a href="https://apps.ubuntu.com/cat/applications/empathy" title="https://apps.ubuntu.com/cat/applications/empathy">installera</a></span> det från Ubuntus paketförråd. Starta <span class="app">Empathy Snabbmeddelanden</span> från <span class="link"><a href="unity-dash-intro.html" title="Hitta program, filer, musik med mera med Snabbstartspanelen">Snabbstartspanelen</a></span>, <span class="link"><a href="unity-launcher-intro.html" title="Använda programstartaren">Programstartaren</a></span> eller välj <span class="gui">Empathy</span> från <span class="link"><a href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen">Meddelandemenyn</a></span>.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Du kan ändra din snabbmeddelandestatus (Tillgänglig, Borta, Upptagen, osv.) från <span class="link"><a href="unity-menubar-intro.html" title="Hantera program &amp; inställningar via menypanelen">Meddelandemenyn</a></span>.</p></div></div></div></div>
<p class="p">För att lära dig mer om Empathy, se <span class="link"><a href="https://help.gnome.org/users/empathy/stable/" title="https://help.gnome.org/users/empathy/stable/">Empathys handbok</a></span>.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-chat.html" title="Chatt &amp; sociala medier">Chatt &amp; sociala medier</a><span class="desc"> — <span class="link"><a href="net-chat-empathy.html" title="Snabbmeddelanden på Ubuntu">Chatta över ett godtyckligt nätverk med <span class="app">Empathy</span></a></span>, <span class="link"><a href="net-chat-video.html" title="Videosamtal">för videosamtal</a></span>, <span class="link"><a href="net-chat-skype.html" title="Hur använder jag Skype på Ubuntu?">installera skype</a></span>, <span class="link"><a href="net-chat-social.html" title="Sociala nätverk från skrivbordet">sociala nätverksprogram</a></span></span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-chat-video.html" title="Videosamtal">Videosamtal</a><span class="desc"> — Vilka program kan jag använda för videosamtal?</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
