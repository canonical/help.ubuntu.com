�PNG

   IHDR  G   �   {��   �zTXtRaw profile type exif  xڍQ[� ��;$��@�n���@P�I���!����=����KҔ<BT�*@�3�����#${2�ƻv�!��y�J�����j��տ-*P�>�j|���R�d
8̛�nl�)�Yo�(iɷ�훿G��p�SȂ,�sN
\N�Ͻm�RM��^�Mt��"����b��{v���ȁ�0��WB��|�S����\����ޚ�v���  �iCCPICC profile  x�}�=H�@�_SKE*q�P��"��
E�j�VL.��&-I����Zp�c���⬫�� ~���8)�H��K
-b<8�ǻ{��w�Ь0���a��dB��V��+����
�js������G��w1����ѯ�-$�8��6��̦]�O,����O�tA�G���q.�,�L�̤�Eb���j���OG5ݠ|!��y��^���=�#yce��4G��"� C��:ʨ�F�V�i�O��G\�L.�\e0r,�
������Z��I/)� B/��1�w�V�q���u��+��6��O�-zl�M�.w�᧚b*��)
��}S��ּ���8} 2�U�88Ƌ���������=���t�r����  \iTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:7abe2e2f-dfae-497a-be43-f4ce58424079"
   xmpMM:InstanceID="xmp.iid:bb8ad924-dcb1-4a6f-8cf1-8b1f10eb7fb7"
   xmpMM:OriginalDocumentID="xmp.did:caa19f0c-47c1-4726-bf90-f5ed59d4bb83"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679602035973940"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T21:07:15+01:00"
   xmp:ModifyDate="2023:03:23T21:07:15+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:be986261-ba60-47cd-a405-150fb54a2aa8"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T14:56:59+01:00"/>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:0e6b05d2-127c-400c-bac3-69319d337738"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T21:07:15+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>K���   	pHYs  �  ��+   tIME�	F��   tEXtComment Created with GIMPW�    IDATx��i�]�u.���g���*UQ�A�(N�,K�,Q�,8"I�-Iڱ�	�F����0�h���� � ψ���a�ىӖ#�,�e�iI&)��HYs՝�ޫ�3޺uY,�\�� V�:��3���5/ܱc�������h۶��q#\�R��=��<���V30X'|�J�R��޲.\3�RJJY�Vk���6�jkB�B�`��Ƥs}����j���I#�	&�f��`�v�Xܘ�6��vvvZ��n��AX�U(�"�D�\Nan��a5�5%�Df��������,������u�8�x≭[�V�����/����y�7o~���8��dN�8���~����K}����c�}�#������_~ r�������z�+W�|��_?u����|�������?��ٳg�mz�}�=�裷�z�K�������k-��u�Z��h4��V30X�I�s�#�t�����;::�\�r�m���_������o�}�m�:t��ٳB�Ç�ů}�k���Kw�;w����>�{��T*�7
!z{{����N�ј��(�J���i�z������z�ڵk����?��g>�s�ν�曃�����s}�¶m��o`X��`m@�&�V�T����̙3R�{�����=����[o���+���j�Z�/�˝���B!d����|>_�V������+W���;;;'''ϟ?�y���@WW�eYSSS�Ν��j�\n۶m�������r���B<���z�駟~����D�8���������rYot��'�,������<��f�����/]�ڣ�B�����=��7�񍙙���"۶�ժa5�jk a]�\8y���Z�6�d�z=�J�q�CCC���������xx��?�я~�ʕ+===�m���;�|~hh�T*}��x�7>��tww�� ���w~��oٲ�K_��իW�o���jR�������>444��v����O���?~���<��#���G�UJ9r�u�g�}������������k׮:t����ԩSǏo�c�,˄���V�ϒ�8Ξ={2�Lڴiӧ?��;w*��]���
]]]_��ט�ӟ��֭[����W��/��w�}�o��o}K����9r��?��6�^y�g�}vttt�	�ܨ�z������wܱcǎ��z��_���s��կ6�Z�v��?����{�-��G������|�#W�\|��G�����_ls���V30X3���v�m����ӟ^�xQo�x��W��͛7�ɟ�ɧ>��.?~<ܿ�h������۾}��3g���Ξ=���t�ꩧ�ڵkWwww�l4ǎ;q����|bb�������?��c����8p��Ym���Ç���k���o⬦	��?��ѣG-���7�y��w;v,��V30X�`f�Ts���/���{G���j��R�Vϝ;�/��/�7�����p)e�Ҵ������|��ɓ�W�������^8������eY�T�uݯ~��������ww�����{��a۶�������>q�D�^/���z�V�]�t�q!�\����200�f`�2�]}��gϞ/|��B��g����*
o����m�n����W�
!���x\�=:;;]ם���������Q���۶m�,k˖-�w�>y�d�X|衇�i|��?{���8:rdd�_��_���{�<x�?��믿>11q���C�MNN:�����_��_��v���H)=�kS��{��{CCC�Z����9299��/~�������f�DT.�����-L*�..\�p�ر|����DԆN�ػw�SO=��ё�d�9r�=�|�K_�f�����,�\.���>q�D�\����{)��Ȉ��j�}�^y����!���o=�����g���g����~����a5�u 4SC62�L6��+��y��>L��ŋS�T�P�I��jurr�^�����B������q����ԦM��Rccc�\�P(hB�m�ҥK��������T*������:;;CO������Bttt�ӫ���ӈ#���ő����X,f2���䤮r��P����'�V30XyQGG�i��juzz��j��M7��`�@)U.�MN�lx�W�T�V30X{I�T2����T*����c��M)��f�+ ���̌�4�jk̬��g��T*�a{D)�*�J�R1���a5����OOO�J%�qtm�F��KѕR���V30Xo�V�Vu#c���-b`````X���������������a5�j���V3000000�f``````X�����������������ဈ��R)۶7HW_�8���F�Q�V����jX�`���"�ɤ�i�d�]�m۶�L&#��V��J��<Co����c��t:��d��!��f��t�T*U�U���=1�f��a�v>�wg�N�40h"��r��LOO���k�i�[��U�b�躮�4�6@D�u�Ţ���j�W���m��
�����.�7�f�Ju�b�hY��l`p�,�P(߆a5�U�T*庮�xw�鴹��V��t�� "�R)`[�ֶ�����3����q����߿?��^�z��W^9~��I3���mRJs+֞N���e�º�4��~D�]�v=��S;v���J%��8p��[o}�����<��uݎ��b�����F>��m�5�����m>6��tvv�R�z����=������J������t<��;::t���)f�P/��Ҩw��V�C"��\7O����S��3��'?�я~�����ɓ�z}�޽������|q�u<�{��[o�u˖-�B��ŋ�ڴi�����:�'����mCi>��m�����1<<|�wvww��������ŋ+����Ɩ-[���&&& ������oll���D�����[��y����V���������k׌tm0�駵a<��S͜O���ޛ��=z��q�i�z����?��<�{���_�����?44t�����I۶S��|�6�>����6�\GG��O?].��������R�Z�瞛������s��T*��{��֭[O�:�f�ԫ��Z��j�����R�d$j�j�&2mX�`���|
n80::z�ԩ8�j��_~��ܹs�|X-��#����h4��r�4�nݺgϞ^x����'O�ܷo�ٳg_z���/���eY;v�x��g�FOO�]w���+�LNNvvv>��#[�nݲe�ٳg���
�x�������<��{ｷ�����^xA�Kx��͛7OMM=��s�ϟߵk�}��g���M�N�>��~�X,����O~�w�} ,˺����nf~��_x� ���<x�`.��կ~511ڬB��z��_~���{��[o�R���K��կ��V30�f���6������l[dtts��|���<��O<��/^�t��h��|>�СcǎMNNvtt<��CO?���K�<����pgdd��vG�"�j5 ����~��U������z��^���>v�Сg�}�X,~����~�=��������:11q�w>|�����ɓ'�;�J��=�����o��������s�=����Y�Tt$r�֭<���~��j�z��f��/~���={n�����R����;vlpp�S��ԥK��xS�&��btt�u�B�д�����'''��!������7�]�v���'�|r߾}�����>��O�:u��ɓz����ɓ333!퍍�����ܹӲ������ѐ������ڵӧO������?���.� ��sϽ��;����^�vmxx�q�s��1�ޭ=ǩ������K�.���л�{���+W����ؼys6��-[��ݻ��_,�J��:u
�]�6==���g�i]j��&[�`U`����_�СC�w���/:����>�!)e�F������g�y旿��;>���\��������>�W���������w�}�ԩ|>���Y�"�d2a3�j�Z��t�BS v�ܩ��J���J�/_>y��@�:u���N���luTO�-���*�&''�Y�=ϫ��RJ�`i#�G�V3X�'����^���?����\����#G��߿�\.�={�������W_}�\.k���˗_~��C��7�Μ9�iӦ��^�u[f�$=s  l���
�e�ڵ�^�������z<�g�&��j���/~򓟜>}����6�:::4���+�Ԅz���J�r��۶���o����Ǐ����4j�V3X��8�D�����}�{�J�����������g��~PJ���~�~KI{l۶�������z衇R���˗��_|��h�{�m�����ɓ'}�����z���Z�\������g�ك����L�df"���K�Rw�qGgg��>55�e˖\.GD333[�n���aۈ|>�m�6=4�q�Z�v����o�}۶m]]]w�u���&ȉ��cǎ�q����J���ή���[���z����Z��W[�Н������[o�U*�l��<��<��ѣGo��]�v�R����}!��8۷o���{8��:z����D___�Z�p�����w�166���{��ŰPl�Ν�Ν���SSS{��y����U6�-
�Ν�RNOO����{���{�3g^z�%)�֭[�^�:22��fff�m�v���3����+WJ��իW�l�r�=�����>}�������/���4���z��|������~��:�W�V?���ݻ��w�y�7�R;w�<��.��>��+����
�K�.�l���z�^�V��9��;�]X�f�:�~a�g2�O|��v�:v��3�<czjl@����t�\6���`�E�'���r�ch����O?-�ܶm�eY��6�������V�sE,
�L�f>!�ɸ�;>>n�m���r�<55e$��j��\*�\�]�4�	�_���4�J����5
��n�y^�����`�������V3X�(��F�40�!J+�J74�`��x �9����fM���PJ��a5���{J)����ʹ�3�8�655e
���F���\.�#�o��f��9���g�FCOS2wð���A��w�u]۶��Xoq�3g�F5?��S��6�Ű���xok�Z�^'"˲���m���(�)�<�SJ�5ǰ��5�JK)����p����a5�g�)W�ی-5֖�b�a�ʃ��$�H�j���6#+�������
���#�*A#��m����2��ɷ����0J�jd���h��l��Gv��h3Oy��h�L7hz:+Bo�J]�2���b=����b�tx�FT�S�Yfn3�V�V(⾬�6�l��9#��_�.�݌L_W ��,�;�����ڈĪ���l��(��[�zYzk��-`�3���_��<ӥp@�f�j���Ik9�����ň��X��et��b7b[�6c$ae�cv����թ�.�<�"[�����������q)�-�M�5��.�+�H�*Qɗ��>��{4s1����?�����r�$�ץ��,|7�N�Em5Xi-�/��(�ވĲYi�ܾԄ���v3�fdt�/g��m�Ķ`7����7�����<�dTި<�Xqy�y�-�Y�v�헤�|f�t�9��Y�� ���_&���*��-u�9/�����J��|9KJl+��?�Ϯ+�F.WV���n�s{n�0��K�r��u�n��&�� ��8x�H,���ߐ/g�m�X��\�Ǟ�` ��̊X��
X1���"	 KV�� T0+I1230+}�bŞT  |���� ѽD�� Y��7`@��?#D?���F�� �9vg8�b f`=$#����oA`��	�g``����'�w�!�'���s���Ե������4�f�R��2�D��_j��5��7���g阏HyX����#6ky�BK���ƒ����ߨX3HF�EĊ�=f�+Ќ��b� J�b�XzRs�� ��` D��_��  	�S  �Ei �@���_��� ⟀MO.�3iּg5#0�Z|# +�*#����1�,��/����H�|i�qP��k�W���\���.@�1"���0�v_fb���R�/�J�I��R�y�G��%l&f�m2��	�}`�9�O���1a�`Hiz�G��;)���@ 
6F���1�}ڣY��~�7�:���Մ7�9�R1Қ������sX"J�ml����6��4�7�����;������������?0����&m��@_5�[���bb�`K�`l��pǔ�)dI�:z�0K`֥5�qY���4�V�z#b�~0���{���O2���|�gǑ����W/}�� �.$�!����͒��0�<��9�!��V���=�H$��Y��_h!*M�"���V��y[�θ�I�n��۲f�7�W��� *0200\���#H 1��}��[d���1�s�S���7�c���~p��C��F���SZDc�شC)�K..��0!�&oP��|��/dl}o�=��5q[Y�m��.�so�?rC��ԇP)W���	�d��@�I�C�f�Z����@��A�TJJ[��Wm�{��Sc��HS�$���[B4E��Ȭ�"H:����˃�A��|�{�NZ�ɍ�-�m����Y|�H^���c7��\WjC��{��_|ň��d��Q:`��rH荬���c��Y���I�w��
Y�㡊��^����Pb�@lR�)�ȴR@B�Ů#�6XB9��D
��s��r�1�N��ܒ_o
}g^�F�F�U�j�	�ˈo]O��V�"@�&�3����5�U�X�x��O1��H��c��X���j	#D�\���"q��E��������D����&�e-�Z���q�%��Ad�S�o��e"����Z;��l��w���62�-��� +:���N�֠x�G�/+��!�B.MDU1�9#��x�5.ƈ��,�z!Dk6��Wy��3K[i9-�v��sj�%�m�5�1����R�u5V�萰��#��9&�
&-�l����g�,pLs��!����bڏ�&T��D����G/l��5	��Ϥ1QZ�*<kZ
GN��pS��
��|�p���WH��Ji�Y	$	3+��R��p���kVD���bZ��]�>�1���(Ü��i���ۈ}��(N��@��C�6��pp�C�U)ftp����M���u�G�8�"3n���M�#M�,���j�m9�����*'�o� LYIP�鬔o�+H�h�����DI�,F=v�|2Ǖ���
�,��S�#�f�~FP�SG*
c�G[8.��	-����p���ƴ�9���K�$���
��X�b2X8�A
�>�1�R*�r�w��3B�I�u�cfh
��pDW���o!_!�$���3��S����D�!�8Ę9)����P/��Z���`�e�_?f�[�>QiJӏJ:��I�_Q���EJ)�2:������ ���: ��I3F�&t��[l�>Z��S�SZ�r�bst�S���Q�"�0��}9*r4)N���y.����T�����k0G� Iދl��Ozl��w��V&��E�������0!�.���_�	=!m��΁�T�^������:�b�C<����y�r����Bi-q�c��k�k
�l�����MI�C�0g��)aY�J�L3?�����(�t���cD���4�눑_'.:�,��CR�	TJ� 5���0�'�23|~�E߃d�d�5410І����/kOl��s���8a��R��TJ�A��`Z�f -���0�O'~?��5d&_�d`V $���S�%���3^,}���T�`5��0���8�VvO(,=ȱD
�X�U���ǘ��ܑ3!�$�p����������Is�op�RJ5^$'*����Q�����&��0��9饆X�|�(z��g�bL�n�8F.    IDATp��eɜ��ل��K7�J�>�$�$,�D>�
w�8����x8������2U1o�p�M֏ba�'�^���S����w"�&��		?Rq�%#�	ߥ�gB�l�� �y�a�8��^G����S\7>0+�)�vq��1��7�	SfE�xiX`�,6kѩ��qIE���-��{衎T�5B⁄Y������1MZ�5%)%R�0eI}<22;��_�y���&�	�|<�Is22ƭ�Z�|��gw�����?��X��[��R�n����DIa�\2�B`���R̺����D�0R���:�V2�b`Ƥ�b�3�-r�0f���\pEai#j}%���,�V�!̱�` ɱ�?G�A{b9VȨ�������C�n�s�Z�z��hJ�Q���@H61*�4�� 1����&�FHk:4��pqB8�'F����i�-	�&��R,�������Y����v7�GI"�� N�D̉+'v<k�\Bn��s�y�[�*�v�R��ܐ��wߧ���k�� �%�Rjzz N�ZǯX���j��	!r��R���R)eY�#w����]�F@\�u-���e��W
d *���A�E$���@�&��(�1��^�|J�\����
?q(ʵ�1;d��xđ!��h'����^��3T��L��y���Ĉ�d��|�3ǣJ*t=!H�	�ќ4,"�^]ro�\���WU�b�Ɉ�bҞ?��b� gH&��RG�"`�'q�3C�q����"�f@�P��B�,V�JA�t�졦l����Z�@*f?���5?My�Q�#Ni���NŊ�u�Z�i��$�-��\���Su����ٳW�\ټy�mۖ�r��?��χ��6m�466f�vGG�bzz���٬5�k���{�W*������BM�Ν�m����ƺ������y���ěgĩR��������b���oB)����U��������r9f�z�������@:�r-�H�Pc����PZP�$H	���=��_JŗD d
|U*Н9$F.1xґ�����ci���)�~'��� ��sC�|F���1E�/-��zR��������3��h@��CJC���=%���DI�K�n�c��O��m̂}-'�|G �(b.GPJ)���vO���;UcP����
�cTՁ1WQ�6D Nf�rC4�QR� Y:�Hk.�����8�>��O���D��d�Djt��j���dZ�l�e�g�ߐ��H��j�R�l޼9��,�!533s������}�C����8��éTʶm!D�T:r�H�!�z}tt�T*�j�_��F���grr�Z����k}}}��i��Bhsmbbbo��[����į~�+DB�����u˲�(�N_�p�X,�v�m[�n]��?w�\gg�6K����H__�R�e-���_�8�4�ؓ�������&[��c��vB�?7����o }[���~�_ȭ���l���<�-��������R)M�M���2�ګ5��D�5$��o��N����Ź!j� ��~>i�I4�Cn�F@�Qz#47�8� �4����:��jnU��I��F����m�[��o�Y�Sop�a͵���m�i5<�4*�J]]]��j�b����Dt�}������D
s���ݻ��B�СC��+����#UTS"ڶ=00 �L�R��<xP��eY;w�3������[���]tl۶m˖-�m�/���K�R��{���V�[�k�B��o��/���gf��K�R�T�Չ�I۶S����q�U�n�-WʩT�V��/��SSS���qa`扉	�u�AD����r��h�r9�<�Άށ��[���S�2��h��ᆺ�7�� �B��-� 1��+>�}�Oѕ����Af>ikM�Ta�Oh�(V�~gX��݂PjZ�X~�dHQZ�x�d%~�F�z�6�`g9�ÝcIѱ�k��P�khj:������*���F=����l6��.�ە���{1���bӦM�g�u��?���x����{���?���¶mMi�TJW���P�Q�����z�5��� �� 4D��T*�%>�����g���yf�p�BGG����=�������.]�<=222==](���_���۹sg��8z������#�S����|�X,V��7�x#���۷� V߂����]�x��뺡��o<�S��]�H� Q(L��x�u��C �K����	u6��e�����Laa����aM鎔LwA\M�Ńm�`k@f�D�R�O����:��y��ԒVl��Ï�%��q+� ��G�'l�¶�\&Z�-ef�vr���4։�|��<�<.���A7����8+@&���jZM!"!DOO�m��z}E� �˅�������Q���'OD���+��m���O|�z�;v�=�ٹs�"�Wa������6��k6�ј}C1�da��3�,��FyA�~X��3a�ć�Q?��u�?�
ىAaH+5��@�xs�`��ȄN����W�*V  A���hץ�Q�%���do�d�D	&��l���DԖ�p�-Kd���|5�]L��DԴ6,'�h���7��P���b+�X�yq9	ݼ�@[V:���{B�X[bppP_��Gg�O�H��t��\.�ٲ���~���>�/�Y�Ul�Is��bP�DR)��B�b%��������q�� ��DD:Ñdȕ�X�T�����D�������̲�g[� P�jh��iPtѓ\�:�'h=�'F?�NSM��f�Q�!2J�(�;���~�DX�>���'��6X�h3ci�b� �R�� �%��|��n����NY���=2V���糸�MI��I�����#;�E�O�Ѿ}�]�(��Q!#���Y71R ��<�`������+��\��4?ݑ�b3BM�X�P#�i <EAkI��9�We���w��)�Uܜ��+���f!����D[0�Y�%�965X�|6�:}H��B�X9����{��5�dq�NPG΀��i|������y-&aИO@��Q�$1
�(��&�a���&���E����~5�+�Qw+!@�Qw5���X!GT��@�����  �KnH���'��Sb8�C) ����RyjV-���̳��&(-Q�����3���Q�Ơ_�fk[͝�e��������СC�J���CJ)��9�a��eYRJ��:�|�V��;��z�V�</��\�vm���MI��mh�����{MOO������U*�T*�N�-i���s�zz�T��3��)�u�h��`p���\�x/jj�9�P#(�֖���&	�C�/�W�R*�gf�[P���uSXdn�ɠcia򈅘�@ �M,�S�P 1X��аEP���.��Y��L�� �ܿ8��x��[��b^�����FrK�[�Ͳ�Q�%���F������Y��o߾'NT��L&���'''������Ο??22��㏟?�P(\�xq���?��-�r�ʕ+��mڴ��;�ܱc�YE��j��Қ'�c���h4*�������Ի� 333������۶m�����B/��7�Q�~AG����#�V�ͳ�cV�^�އ���Z�(<d��'�3�`D�x$""��,$"$B��@/��JI� ����|��ͧ1�;�c�Я��ZH��)�/�T��B���g�$K�
��Rc��]�-SU��n��qY��� �RN�#�q��ț�7.��v�e`)�����#G�hSlfff˖-�L�V�U*���N��B7�pg���ڹ.���'?��ﺛ�N�3��t���,�x�;�tvv�R�T*��ӳ}���=m�����/�T=	�~p(��~� �ʐk��(O�ꯝ�)���k��O��	7�IP룎���q�N��v����aa�E���� ���y���5O��ou�a�%ps^�U���6���|�OQ�ˠG0	�%Av75׹D�m2"!4�	H�"�D���.��e�,�EĠ��:κ��R� I7΂��:�w�ʠ�+FɖBK����Ƥ(Q*P� �6O�u�R�<a�Ҵhhܗ��`���ϖ�+�{��,�;.�!�eY�
-�Ur',P�Ю�8o��@ˊ��|֬�B���G�.]�����M�_�Ul~��ʦ<9����ޕ>�==������3?:Q�:6��Y�ʐ��Bȧ��e��p�V��7f^8Ӱ	]�w[�4ZB`Υ?�?wK�������V[`Ɓ��V.�#C�w��|(ߙ�V�$��Cd>"��ȴd�+!
�e��=��G�u5�H$I�"QZBؖ �<�@�(�"F���S���H@B�����k@B H�2����,XG�t�ʠI3x��@[`ʂR=���z�yJ���O+]}?�"���h�u�Z�%����ҟ�Z"��&��zn�̌.̒R�ਸ਼�u�Hf��(26v�c�%�'��d	�rMʖ��]��E6�%�;���d	 �x�\H��0ȧp�K!�;��9�8ms�� �[	 Ӑv����l
� �W��|��y����������6�$���t��
��#��:5�	K؂l"� �cf�(��0��"/��>���;����&Y�s�%lhx�KU�$H�DX� ��@t,�P\i�J	�J񬒍�����jb��VRp�����jJ��gu5�U�m�X���mW�����?�����FGG���y�TJ{����|^�,���@�m�]j� �=�Y��@�\̶Y��w�D`	��b"�	������)fY�k���B����(A��m�""Į��Xe	v���l�P�U0Ɯ�զ�D���P	�����U�=�A@�m��Q��l[lKv�em�����
+"����-�W�O�Q��X�F�,�4Z���"�)`$�L
X1*Ũ#g��&O@�������'C��J��,�	�h^л�]��
�&�'A��jaG|����X}��ɥ�5m�,�cz���Μ�Y*�(R�������x��udtbb��hlڴ��<f�T*�\.�N/���.��^.�А|�AyΣ,L�(�sE^��6��[�-@&�+[
S��Gfd_Z�X&�sJ9����ީ��6���$,��]|)X1{*�:�}�g�%+7,B����A�,z �ы(dK{Q)�<�g�Ḡ;�p���c6��	O{Z� ��%�@A B�Hz*�@ib��S�p8(D D���SP���˝�҂�p���+���`�![d9n��L�;�ϼ�^�C;�Oޝ��X��6���z�붮P��~�======s}�w�Ζ��MK����n�58�µi�-b�9!�B�#�#{�__lL��-](����X3�6���Lse�[��>:;"�u��`��V��`ǃE�Qɦ�a�Q̓�@�����~���'*�
P��(b��w�eSJ|4b���h�� 5���B�����O "E��m��rl­_���+�(U�:������N�H��J�,GS��S��x��_oW�M��|ꃹ|ڪT*:0�oh��H��###�F�����r�\�P`�z�ND���\�u]��*�J�B��h8�cY�vNMM
������N��IJY,۟��y�j��*�f�W4/p*9M
xff��Y�7�u�Lfv"!b!�m��$b!`.~Bو���+��	���q!�peBVj��=y��Q �� ��bڅ��杠U6YX�Ҝ[�j���x�qX�̱������`��f!�AJe)`b��Bm�x��b�|��ҖO�[0�u���{AF"(`�+�FUx)hY0#�r���X*f��d�@�0e�T�r<�!Y��
�3,�YKt�sB��l�0:����ʯ_�R*�J�ɼ=,������y%��ӧ=�������gΜ���l4�|~xx8�ˍ��y���󼙙  ���)D������4�uk�������t:]�ՔRw�uW��RV��r��W�F�!����^y�h=�	y~M�c�qf=����߱c���hh�Y�.�l�jB� �Թ!Ywd� ��?� =|��l
��@���X�H���2`[,�h���r�Z��δo��l�D���s�b�X��A�b�:C_*�*�Eg�``TD�9��*��%+�Ak��pc�sC姖00"204$#yQ�v�,��˱��j��s��z̈́��QR�bf$Dߛ��5yh7���
l��b^��>6ݸ0�I[{S�-%������Gv�;o��y�z���!F����ڵk�^�v{zzf[ccc���̙3�|����'�F*�ڿ��'J����������n$ߣ�{8�/� )�˗/_������ =oQN	�`K�-�V�-+�����,� !��x4g�"��P� oÞ,� �`	hCPD�B$��.�T�>A��\4���/�\k����˻R��Y*�
Q
��Jb�T�T�S7�7RύP�!Ɖ1i~�?�ғЁ��8�A@�;ia�*Y)&������-����7�(�d  ���3u�dn�2k[�Vښd����R�������?}�j�]�z�T�� �֟���ۈ�%ڶ��f��8�����n���͛[�i�}I���������hd2�T*����̶mW�US	�-׾����.�u8p�8�Y�pQa|�""�M��VL,7g�f������d�Ϲs�wxK��a�u�ʳ%�+�����A���B�m!r뼯��3�*�7Έ� 3 2�z�Q��b	�����C�:�VH`�Š	~�-�Y>���5�  �#aC�Mz'&	�ҧǰ5�N���%()��,t�& JЩ���hgl.�9�	��W�`؍�j�"cm�`[�w�%�}��JRi��k=��WG�t�w=�Ĳ�L���Mƹ��0t���R��� ��lX�v�����[��[�ol� �֛��7z�m��gb<0ԹA�����%ܒ�� T�����Q1KV��I��*���j~��4� ,[���d>��hX��Ր@�U	���u�B��ђ��3H���D���aX_�i�"r-Ym���3ep���_���H9D��#h䕳������6�
�O�B,]ˌ�
��( �8��������А�yJ�T*EDVG�
�MNN�����i�u��b��W��������N����t�^wGG��T�R׮]�V��\�����tZ�.�SJ�	�j����z���ק3�2����湩�i�f�*�1>���I�@��&� 
��* "�a�c�� ��*�Gm�?��D���*��ف��,�[G2�T }CBffɬT4h���
$(�@ظ���&VBּ��
nX�lU��R˓�O���t߳�˸�%�x��6�j�q,����R�t��Ł���'OV*����J�R(�m۶��\�ծ^�JD:�5C:��333###��w��H���뒙y||�����|����T*)��F�\޴i����۰��-���ԗ�cǎ5�j7��-��ܢ��y+�[:~������Q2F���#u��܆�"
6!	Ҋ�b'h)�#٢Ӑz������#��e�.�D��0/%D��i��������T�5LF�5�lKQ�f����؂0��a��ђRn���T[.�۲e�eYCCC�FC)�N������{{{�
��D>�߿��Z�w�޽{w��j�B�:��L&�}��Eo����d�&����0�̇��t�=1*���Â�(*��$d��P�۲,T�89!@f�
Pg�0��i͌��"C@"#&fUKf�ʓP��$�Jq��X�TJ!1�#XJ��tGc��k��V���V����8�&�./��r�\b��\׽�q���:k�����Һ�^�u�`P�2M�cJi7b4u̟�Ċ��*���d���v,�l"���o0� J�Y!���>Š@I��=�1j��1��ŬM= dR)DB@����t���*a5h�LX�˳�u�jn	cnR@���q����� ވ>Nc�����9�]�gx�Ӯ�����.�SA�b���w�B���(C�T*QS�{m�4���c����e�6{���L�Z����\�H0*��V�~���7k���7  ����r�ʶm���}۶��8ж     IDAT�����_�y```�����s�gީJ	�Y����|ʯ��eb?x��n�g�� xK�>vg�ƜA�mm[{���M�35Ax[��[{2���vG)���__n�{�����£l�igcH;s��1�M�|w�]#>H������p����02�Eia�`����Q箰�d���gR����C�c8{V7,�b�x�Q�1�V��f`p����4�a�캮�䢔�z��իW{{{�����׷�o�{��3��<^������#�&�,�8����#��-�5�g��?�u��X��[�-�XL�g>�����5��}���w������Ml�G��8�٢�����|i�j	l�??]u�i[�M�)3�_����Y�\ F@R��;bM�(�pP+`dB��D�d��_Ϥ�?��1`�H�-E�z��1>�:�C�)���f2XiZ��o�haAB��k���_�m֊U�jl��ד����b�X(qϞ=K�J̻`�,��[�!@�J9J1�V�՜�QC���֔L�j�Th]7�
��"ؾ	����RLU-Y\�.Xl��n���ML�T�]�XU�w��G'~���~�,���G
M.�	 ���5�A�6�"���h:HA�!j2�0?E���y�J��mq��ا@��*��A�o��4M?��:}fa�X�-��eh��z��쇥�*��^��}K� �l#X��|k���۵	Ķ��T6p&���M�־DAp`��S�%�cA�E!��m,�s�9�!|hGJ��=��.,,��u�� �C%���������pBb���#'��賟C_�	;#:$��s���tQ̠��CmbI�A3]��t��L89�b��&���c7�`�YC��<�vb��"��###����J%��ׯ�.��0�Bڡl�1 ��Hǆ��)s�)&��K�����&y���)�e���.��x,΍�B�;sH��)��U=D����6�����]9�ݍ�!͑0h1�5v1�2a���Եҡ�!�� ��;WX�oU�[�s��(�<)��%�9ix��Ȼ�����~�-6M&Q��7쟂��1��j��b���� �֢	2�Vbc�j333o�����Ϝ9S��5���i)��ؘ�бw��'��?���qd����nR�|zX��|eBm題���\�?*o��	��%�%���>CA�1���P���\�)�h�^�¢g�� �#�*f@�A� Bd����&��- 0(dLY�@a�,��;�!���<����ld V
�ҹ�A3ͱ&Zt	IJ;~%�������7�͓X�+�c�ǡ�E��B���t����K��{���z1)������t:���,��u+}8=,��z��G�?��4���צ� ��ĵ6GY���2.�%� a��� B� θ0S�l
<�a��'�"�kYi{)���w�;}K�[�T���E�د1�oѡ����lK8d������[+溔)9��k������0n `w!WH�/�����	B����*��d�*"�)�!\�*�UP����q�Q�Э�1jF8ʩ�,+��C����m�R�����l�siD�����p�WWs�^��gU�|mZ�������Q8U��<O������n�q6�{�xI]�T�Ǉ�@W��l!\۶��Fm�\;A�)�$0ى�:l��/F���!��BltF�Z(t�*�(mY~�,��X���${J6<O�	#O!+m�q���@i�w�����ѩ�;��:6=�ܛo5��$.�[�~��ψȵmǲ��5Msū���m��±,K��"?Q�KS!
�1s�\�ݨugY?�l��D���ݷ�� JĂ��=,���jN�〞��s�<��<➂?)����]�Y؂7�`R$b�<�R��mY�%,a�لK���A�cs(-�L��q��8+$\��Qz�[HBw�@��l���(�_��P��Ɇ�J��}�G����1�
�ܖ���-�[7�<�گ<)�T��ɏ���[���l�q�t����ȶ,ǲiW�ZN�VvQ:p��ڃ%Dʶu���불oX�V�ccc�/_޵kׅ�T<�~lj��P�#v��m#�~����ȸ8�|���VW
���o(H]��棅�����Qˣ:��\N��}���0��
��Yg��h�ȱm[���Ү��� �ڡ;����&>%�$��e�t
�� ۱� `����j(U�<ϓ�r8��?+Ś�8JQ� i$*���-�L��X!��{��o����|�5����e[�βY��_Y[MV���֔ˑȍ-dQ ��G��Ar?"�Ix�b1���y4�U�C���Myw.�t����"��QD8Йnc�u��{�7zԒ��c�N0��c��q�3?�0���S�2�)�?�O&����c���{<Rڶ\��-C��c�ֽ��4A	֌>`��S���%Q��~;��� �z���c���(��~�N���JnDD��u��ϒ��2^�Jw�Z}��A{����:69���̗�R�Y�ZWWWWW ���,� �ժN�DD)e.�kO�����L&S�T�����םS�V=�ӓM����̜J��|��S�R�V��TJ�YΙ���m� ��%��q�dȡ!?iK��Þ#1Wd�^1����� l"�)��:�.����Wiԙ���K�����8G��E�g��zR����l:���5V*�b�s[����ض� %�*g/��3�櫘A�e"@`�(��\���a�s�gff���5a�j�={�X�XPJ]�padd$��4��;w��6�K)+�ʅr�\�Z-�B��o���������q ���߼y�2�WCDK�mY�3
D��,����?�3a�i�IC�!���h�O2Ⲩ� ����\�R�=��5�z	#0R�k�L������bL.�AlC�2^X�pelbsg����C���Y�,!la��q��)_с%RwW;�����	ǂm	Ꮬ\�6�-��-9�%߇������B�P*�ǑRj��f��g�������Z�j+j��:;;3�L�eYJ)۶��/���r;v�p]��h�2��0��͛�������2P�%�-�%Ô<�	-�\���ɘ	l#na`��X-���#*$6 B̹n�u���ꍆTL���%�BfMNDL�'���LX���Z�
�>3�͏������b���Ƥ4A��DYgݧ ]��JL�[�E~��@�i��׵-=`>
��S�\5���-rf?6����,Kq�ҥ��˲�����4��An7p���d27�18����������o�R't-+Pk09��1%�!A-#��	����u<�3fB�c`�E]�|�dr��%Dg&[��Z�ו���%+Xr@ DHH�L��43�H�O׹�AP�Ȁ�� �5��4���_&ؖe[>��{�3� ��,�Y+{�Wq�6�˲���z�k�nԐ���/IdX;���"��%
�m���ѡ��o���P�D�iyNU���}M�#ٕ�9�YY]Ruۀ7H�ZH���7�_�������O��;oǀû�5c0�$���Ւ�ԕ�d�{�x�E�F��L�ɬ�@��$3Ɉ���s+�e�P�J~J��nYH}��-�L��뛯cz� 	H�Qb�4�`��=FK{nk?����}�2��v���j�Q H\7d���nV�!�r��d��-���_�WK[b��+;�M�
!�Njʤ��34�M<OH^�9�2rI���7MC���E��}�uMtS�pxO��o�P6��g��a��;FeO�T�f�H3+٩�F�^y�n#��$�ϊ�����}�h��MR���`r�
]�vJzxM�Y<X�C���'�Ыu��Z]K~�lլ�J�Pop�jد���u�:�p{{���~��W1Ʀi��]۶$/�a���|U0k���F�Ri/U�u@��tf��6����kO�"d5��U2Kn��0˴"I��"����H"0�vh̚�@��į?����l]ϯ���Q����:��B�`�{G��������/o៷��L_�ј��&4;i���"S4�����W� I����w_�������7�C�4͇����o��v�^'Ѭ�����5}��02��,*,R�e@Cl�l����.]��dE�8��4��@+��\_[������4�#cch�Ƙ��6fQ�=xG�������Vn�B%����6�yo>��5����+R^�A�˔�U��R������}�8)[$��G����m���߷m�����i���G���׿^��ÃK��B �'I5�Kݬ���:�9�P�Z��1Q>F�q�ɺ��{T~D�&{����d�n���\����Oi7k�G�� zj 5ܕ�`t�,ǰnB�Ύ�C��,�	�=q���<�ݴ��r<��(�-<�m��j�S�Wy�b��~������t����D=����16������if��=��v����ujW͢Uj��S�6k�T�L�����.FA��B��41��T

��sEW�~�Z��Ϣnz���K.ش7�\������b���r��&�f@��(�7:=cEDÉ�㔱��q���r����e{�_�8>ԕ&(3��yt
Z�`Վm@譒<a��	�����ݶ�$��BV��;Yx��o�k�Q[�-�L�@���M�2�8<tT��41^�m?�&�%M�2�6a�4c/FT��V�/�,������}���Ѻy�Q-kF`t{���Q�(����h$QH �q����n۶m��KR����c�v�`�)u�>jaD��pU{'�˕�ݱ�}Ya��B�|n�(�h����"�[��T-W����|S�(��I��W��T���޾}{��Ǳ��^��ݭ�ae����8��g~m�4��j�$:I��XL<W릹�l�ۤ�&����
!E����Ɂ�}�`�m�:rGTqouu��U���#�igi�f�P�G����E5��
�r�V`<��%bq��>|�կ~��_��o���o��W_����ݗ_~���_��ݽ{�����_|���]{P������d��:�R!zP�K_^�#L~�^D������nI�|���>O*t��D�u���4��1�&�5�,Wf�����V�wޮ�Һ��^ $(�u,޲7m'`�W[��qk�,w�L�@�c�����������,�D~�ӟ&���ߓ��/ڶ}�����P����u�%3���8��WF��xy����/�C�νa�.Y��������矿��i��X�U�m�[���ª�&v�I����}���~$�%Z6&�6x���=�?]�����H.������O/���M4_|��r����!������Z�z�#?�b�n�Us�t�wi�lC��Q��IR7��I��ThtO�)I��1Mѵq �)�{������ʋ$kΈ_�7%j�)j�4B����x �1]r��(��vT �v(��b	�n�p[��t^uU�P/��t��J��j�����8�`����uVr�#�:9�-��Z�P�H�S�D�AJ9]m� #D�\o,ܵ�������;�.]$&�f�Iu&_�1r��VZ�N�0�x-^m1����:�V-�����b8{[����TJNw&ɪ�_6;oG^��Ai�6:��ث)�Lu���j8���j#s�%Ner{�G|��#m[ϻcHQ.҄w`��OB�EۺG_Ӷ`���ť]��R�>�&�з"�J�ت��az�ZT�;��,:K���M�,~7o���6	:ؒ��ǖ�\iC��R=��k����9�6�%c�J��6�Y}�m΃pP<���5�-�IY���8&��7�3!�3�_��`c!"V����ʯ���I�SU-�.�Xq8G}"�'�U�k/k~^��r\���iE�`�����΁��vù�S�p�X�i�z�%�8��!��<8�2][IL���m�T�̕�����@�bE�+�#n�Ĵ  
Q��c+����Eaպ�ے�Bh�M܊���E�]1��*T��t �@���H�r��U���f�p�����jKd%��,{!H�Ń����jT���_-��Y@r� �*�D�h�+;&�_��4*/1H���[1}������4N"&�F����;�B��(V}��i�J��$X��"cw��ƫ��@�U�Ɗ�s��b��#�J�Sxx}^m�lWrt3�]PDR%,Ψ�"�J"w�|v5�����V��C�������dO6��(�)]�hT5Dݝ�]ٴ��aq���h^E��E��m�mT�I��B�����1��˪F=���� ��e�x��D��������[�˧jW��cu-�.EȞ&bY�V��Ȯ�v�#gy�RN|��=eiQ���.���hzE�l�Xm�T	�K����؉�4#�<R��q/<ӋIgZ�cf`��4���ǭ���B�<�>wJ���
`Bt��tM����\�BX/�y�օ0�������G����j��b��˱�gBf�r�׵FuҀAV�J��`�@�&	/�)#�@WU���=�j��-��S�i��Мe��f��dԳ.1\F���ێ�)*�=�.h�i;����]ۿLB�������`Y*�>]W��^�kU
3 2X�&�JFc�{�Oq��~Q"��Y��n7(���+OU��w�#TU�S����r��J��Dۓ�[��^D��gi�vmi��z��	'�u�N����Lq$�Q�+�T9�q�!?�~��jL�R����o�;/�'�@�2�Y����_��.B#J9:���x�-`5��<�ݰ{T����z˱�j�\L�?@"GW�*�V<�2��1�S��k;y�D}D���gi� ��Q��M@����ff���|�᫼K�@&l~�i��5<S��t��Ň{�������<��'sH�R�&��!��G�V�.���G�5U�8��sʲ��tT�g���vE!|Q��q)z��(J��:��e�+��a��l��6Z@��͠H�w6�k�`9۩wO�z���!�9io�`8j�x/���f���}�j�D���$�@�����[S��u!! �D�RzԸJ��<��ym�WA]�� QV�32�BN��|�8eD	tFxfV����y�Z�Gy�s[�+�z��
@!q��"y剙�<x�)@�jo�o���7�W��$��8Q��$P����?����c����&rE6��djŲu�x����W�I?�r��o��69�[S55�7���%w�N�L,�����?�!V��� 'A���
�2��S�|�m���gt�G"W!�R���.�Tw�	!(�&��2��9k{5���0�r<�a�F��#t�Q1uݒn7+=��w�nO��f@b����������7��S�P�!��i���)�>hy����HsC=%������?|���Y���Da�h�}K\eB�\d����.妠���`�I!���yb�z��._{v��Ur���
�ꭣb ]�O�����+W*�n	�,r�d�V_���	V��I[��k�94B'�V2/���䎺�9��P��ux�AE`9�#O˓����5M�B5�B��C�U>"B�L��o{��wn��G�p����DN&��
�Vۣxأ]�{r��;$��}��k0L�%�kC�R��
0���1fu(�^�p��ﮩڄ1Y�z�수������u	�H SL�j����؂ɝ�@C��nۃ!: E�gS���:��SU2�VXc0�>ʥ�ȕ1Md�ߡ�{Y�a46T��Vˬ:��|�5�:�vD`����8:� �(s�8#U�g�W۪���X�]8>���������6]A�~�]x����j�p�g�;/�c!<x܎���X���Ʊ�M��w+�EmZE	�ư���@e�[U���XCK�Y�#ɓ[�����9�t8�A�rÃ��u=n��R�,�����Y�G�������7k��J�N��c*E2W�kڈ�����>�\-�9����_���Z&F!-ZK#; r�Q=�[;@Mm��X�czl�%�&���vL�_>�i�S& ����]2Γnr\n��|����궕�7��M��6V��(  IDAT��< �/���@��<NQo:���CbǙ���f2���֟zc�Ie�i<��J��u|�������o����b�~��o���e�W��<��b���j'�.�9�M��eVꐩ&��dd+Y��w�uN�N�[6�M��s����|�B���@#����S7�.�G�3�y][�Z�CV���&�29 �ӱ2l��u�����u�!;�P�)���C�<�g�q��l�mT��q����]�7��eJO�V�����{��/9��^�G�{`�ٶ��{�<M��Y�͕�!�4vb9��9���Jܨ��[�=�`��� c#�r#M�g�5�/_�8����)~�ض�}�iy`@�ְi�����
XQ��1��Q4D�(�I�^}�F���b��y�}WRS��FY�e�E�0td���%?ɻEQ��mD2��ʌ���p�lL [�*�JU:�SӹU~k5�E�������=/[$���o��/��_|����<i�n<S�܇֒�_������ !��*fSz������S	Z�Azi��]ku�7璆��,���'#�r�NG����q�w���ZS늂Z(p$0���ر�d䈞7����Ш��<���37L�aR����6�N&P25���\! �:Јֱum"\\c�lL��!a�����S�>sx8aA���u�+	������W�����!�`7�A���p7s:ѧ�ns	 �pJ)F����?����f�FX@D%�'���wە��3�
�gc�.���������N�q��N�Qv;|���*�D��غZG2d7$���d�5�ĦH�H�k�l.1=&ЩA2B�>����P���K@�M�A��C}[�����af�F�.��4h��$�E���֔l�r�n����q��9��9i�Ə� ��������w��]/׊%����]��8����J�kEr�`h�����V�P��T�Pֆ�X�m����\����<��� <L&�:���M5h�7$�mT�k��A�6-o�b)M����"�F���a�aH���I�qR�0���[�	�I�kҀM��o[�	\��V��!�$�����������e��R}MX���!;����	���\���5U��U9�%ot��F�P+H�qS��@":��:�%�X6�}؀�\仏+?�i�j��b]��������r�ōc=��\֨�r�}�7h�X�.���F��ۦud��@������C��n��sbC4�v޶x��rRu�7�D�M�È`i<M �6m^��~��<����wz�8��@����9:���3�7��uP �l�Yᶱ��(o�j��fѠN��@lw���d���j�C���FĬ	�&j���?��hVWw� X�6JP� Ҙ�tP-�6&h�/�%��Ei�<$�E�siO���#�F�m�m@���Z#ց�˽�C�|h���րh�i%�r�%]��g��h�D�6	������Sk���?{�s���{[Fj�=�#U&�A��FEa��5��K��@�H�%�R��g�E�~��kI��f��ʦ(�Z��;)����Q�V���/q2`�j-��@ ѻ����O�_'vB�3i�c;\L�o"�84"�1O���X���W��α}b�Y��,S�0�.~zmL�[:�G�]��wz��� ��k�Ϛ<��2PIЕ��%��b��dc#ku��S=R�>�]$����6-�՘`T�ȕ�]�S[�4"h+ oݵ�$_����q��$��4tF����m�ۘ/��~L�x\�������u���:����0�rݤ8�~:�9ǯ�0�U�Q�ov���L@T�
p��&��)�>n�RT^��t����>L���e��O�,��v�����/?�<��I=#�	Q���L.ݶ�������&  f��A��~�\��*��f�x8}��I<t�Y%��}��l�6-�Zl]�6?�ț��p���i�ڑ��9G�
�\1�ή^�'4����U��8�2X� �}L���K
ɱ�i,� ��E6��y-!�X��L��� !}�C�}�kR�G�20A�np�b�j=��W��&��'pr�j�1i
Ϲ4��]ܠA��8Z�^B(��Ͱuݵ�D�G0Cc|��l�v�P�p]��:ܯԥ5��~���d��]�H�ĭs:YRAY#��.w�	�@R$�EnEBJ�Ny��1���(ҫ렘ͶW��Y�LS�����0���X ej#nK�&Ѐ7Z��޿�a$��J{i���><H�`�D9�_/]�m���n�:�����LԒ*�2^���L���:Kk����oNA3��j�k��$vv��$6�xQ\7��t$��a��%�ᄟ�	�jњ�B���8��KsӲYe��	4�7��t�f��4��v�R�\b��>�@����ML���k9O�֏���:W���gu0��E�m�6�Y��ar���zg��^<���nl~W�?Wm��؆����M���k���p�>n�v%�4����R�ޤ4����F�I����K��֯��h{�v��y��8ri{�Ns�������~��뫿���a�[���f��H��Jˏ��ē�,Q��qg��ݦ��wn��0d��@!��}�wi+�
�iP��Ƿ��\wo������k�*칻��?� .x�H�ʥ]o�v0'����4���c�_|�)ظ<=�Ԣ���7�μ��u�C��M��(*�}��
���h㐯���c0�Ǩ�����L0>��ܓ��AË���$H\�`����z��r���ح,�^���q|Ш�=��4�b�3GY��g��������&�GF�5$��pr�����c
�4_�K��>D��Kv�Nu�i���L�'�ŞK�o�T��Ƃ��Ab�\?ȷ��xu���v�KI�j�G�G��ff���.$fv�,�)#T<D(�$:��؊�	��]�3Ma7'���,����F%�I����Y���Gfc�m��hTYU����+�׏wiů:6L��G��m1�����Es�Ϲ�����s�l��'䂭����ڑ�l$*\�!{�K{����@��p�,�\^{����-�s%j'	���x|?OdA�Űq�#� �v�cۓ�͑DH</B��0�����j{й�eϘ�=��t$x&�בq�r������\ι��h.��:��6k	ɯ!u;&BP�|O��`����j�s<v��Þ�}�Õ�O��uy��v�K	���#�A˵��J��M�~��c\݂�O	ו��D�5K�]��B�	C��<�=����X"��e�O����&mO�$N�<p����3��~P��ԗ���U}�3g�K��A��仲�$m��?[ �I��Z�ڑ�أ�K���p���j�9��[ q���|�~GN
-�x%x���'�>�ⴰ_D�v���1l����S]�'�a�ħ�k�Վ/.-]�
�����[t�_\N�P��י��T��Cť��l����X�\ҲO��=�7/�X����Vxv��NJ    IEND�B`�