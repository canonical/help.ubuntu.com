<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skärmbilder och skärminspelningar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 25.10</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="tips.html.sv" title="Tips och tricks">Tips och tricks</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Skärmbilder och skärminspelningar</span></h1></div>
<div class="region">
<div class="contents pagewide">
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Fånga hela eller delar av skärmen som en bild</p></li>
<li class="list"><p class="p">Skicka den som en fil eller klistra in den från urklipp</p></li>
<li class="list"><p class="p">Spara ett videoklipp av din skärmaktivitet</p></li>
</ul></div></div></div>
<div class="media media-image"><div class="inner"><img src="figures/screenshot-tool.png" width="500" class="media media-block" alt=""></div></div>
<p class="p">Du kan ta en bild av skärmen (en <span class="em">skärmbild</span>) eller spela in en video av vad som händer på skärmen (en <span class="em">skärminspelning</span>). Detta är användbart om du vill visa någon hur något görs på datorn, till exempel. Skärmbilder och skärminspelningar är normala bild- och videofiler, så du kan e-posta dem och dela dem på nätet.</p>
</div>
<section id="screenshot"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Ta en skärmbild</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Tryck ned <span class="key"><kbd>Print</kbd></span>-tangenten eller tryck på skärmbildsknappen i <span class="gui"><a href="shell-introduction.html.sv#systemmenu" title="Systemmeny">systemmenyn</a></span>.</p></li>
<li class="steps">
<p class="p">Skärmbildsöverlägget ger dig handtag för att markera området att fånga, och <span class="media"><span class="media media-image"><img src="figures/camera-photo-symbolic.svg" class="media media-inline" alt=""></span></span> indikerar skärmbildsläge (stillbilder).</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Klicka på pekarknappen för att inkludera pekaren i skärmbilden.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Klicka och dra området du vill ha för skärmbilden med handtagen eller hårkorspekaren.</p></li>
<li class="steps"><p class="p">För att fånga det markerade området, klicka på den stora runda knappen.</p></li>
<li class="steps"><p class="p">För att fånga hela skärmen, klicka på <span class="gui">Skärm</span> och klicka sedan på den stora runda knappen.</p></li>
<li class="steps"><p class="p">För att fånga ett fönster, klicka på <span class="gui">Fönster</span>. En översikt över alla öppna fönster visas med det aktiva fönstret ikryssat. Klicka för att välja ett fönster och klicka sedan på den stora runda knappen.</p></li>
</ol></div></div></div></div></div>
</div></section><section id="locations"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Var tar de vägen?</span></h2></div>
<div class="region"><div class="contents pagewide"><div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">En skärmbild sparas automatiskt i mappen <span class="file">Bilder/Skärmbilder</span> i din hemmapp med ett filnamn som börjar med <span class="file">Skärmbild</span> och inkluderar datum och tid då den togs.</p></li>
<li class="list"><p class="p">Bilden sparas också i urklipp, så du kan omedelbart klistra in den i ett bildredigeringsprogram eller dela den på sociala medier.</p></li>
<li class="list"><p class="p">En skärminspelning sparas automatiskt i mappen <span class="file">Bilder/Skärminspelningar</span> i din hemmapp med ett filnamn som börjar med <span class="file">Skärminspelning</span> och inkluderar datum och tid då den togs.</p></li>
</ul></div></div></div></div></div>
</div></section><section id="screencast"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Gör en skärminspelning</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Du kan göra en videoinspelning av vad som händer på skärmen:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Tryck ned <span class="key"><kbd>Print</kbd></span>-tangenten eller tryck på skärmbildsknappen i <span class="gui"><a href="shell-introduction.html.sv#systemmenu" title="Systemmeny">systemmenyn</a></span>.</p></li>
<li class="steps">
<p class="p">Klicka på <span class="media"><span class="media media-image"><img src="figures/camera-video-symbolic.svg" class="media media-inline" alt=""></span></span> för att växla till skärminspelningsläge.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Klicka på pekarknappen för att inkludera pekaren i skärminspelningen.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Välj <span class="gui">Markering</span> eller <span class="gui">Skärm</span>. För <span class="gui">Markering</span> kan du klicka och dra området du vill ha för skärminspelningen med handtagen eller hårkorspekaren.</p></li>
<li class="steps">
<p class="p">Klicka på den stora runda röda knappen för att börja spela in vad som finns på skärmen.</p>
<p class="p">En röd indikator visas i det övre högra hörnet av skärmen när inspelningen pågår, och visar antalet sekunder som har förflutit.</p>
</li>
<li class="steps"><p class="p">Klicka när du är klar på den röda indikatorn <span class="media"><span class="media media-image"><img src="figures/topbar-media-record.svg" class="media media-inline" alt=""></span></span> i systemraden.</p></li>
</ol></div></div></div>
</div></div>
</div></section><section id="keyboard-shortcuts"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Tangentbordsgenvägar</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Inuti skärmbildsfunktionen kan du använda dessa tangentbordsgenvägar:</p>
<div class="table"><div class="inner"><div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="key"><kbd>S</kbd></span></p></td>
<td><p class="p">Markera område</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>C</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Fånga skärm</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>W</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Fånga fönster</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>P</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Växla mellan att visa och dölja pekare</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>V</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Växla mellan skärmbild och skärminspelning</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="key"><kbd>Retur</kbd></span></p></td>
<td style="border-top-style: solid;"><p class="p">Fånga, också aktiverat av <span class="key"><kbd>Blanksteg</kbd></span> eller <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>C</kbd></span></span></p></td>
</tr>
</table></div></div></div>
<p class="p">Dessa kortkommandon kan användas för att gå förbi skärmbildsfunktionen:</p>
<div class="table"><div class="inner"><div class="region"><table class="table" style="border-top-style: solid;border-bottom-style: solid;">
<tr>
<td><p class="p"><span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
<td><p class="p">Fånga fönstret som för närvarande har fokus</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Print</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Fånga hela skärmen</p></td>
</tr>
<tr>
<td style="border-top-style: solid;"><p class="p"><span class="keyseq"><span class="key"><kbd>Skift</kbd></span>+<span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>R</kbd></span></span></p></td>
<td style="border-top-style: solid;"><p class="p">Börja spela in en skärminspelning</p></td>
</tr>
</table></div></div></div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="tips.html.sv" title="Tips och tricks">Tips och tricks</a><span class="desc"> — Få ut det mesta ur GNOME med dessa praktiska tips.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
