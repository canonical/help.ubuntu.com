<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>I can't hear any sounds on the computer</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> › <a class="trail" href="hardware.html#problems" title="Vanliga problem">Problem</a> » <a class="trail" href="sound-broken.html" title="Sound problems">Sound problems</a> » </div>
<div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="media.html#sound" title="Grundinställningar ljud">Ljud</a> » <a class="trail" href="sound-broken.html" title="Sound problems">Sound problems</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">I can't hear any sounds on the computer</span></h1></div>
<div class="region">
<div class="contents"><p class="p">If you can't hear any sounds on your computer, for example when you try to
 play music, try these troubleshooting steps to see if you can fix the problem.</p></div>
<div id="mute" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Make sure that the sound is not muted</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Click the <span class="gui">sound menu</span> on the menu bar (it looks like a speaker) and make sure
 that the sound is not muted or turned down.</p>
<p class="p">Some laptops have mute switches or keys on their keyboards—try pressing
 that key to see if it unmutes the sound.</p>
<p class="p">You should also check that you haven't muted the application that you're
 using to play sound (e.g. your music player or movie player). The application
 may have a mute or volume button in its main window, so check that. Also, click
 the sound menu on the menu bar and choose <span class="gui">Sound Settings</span>. When the
 <span class="gui">Sound</span> window appears, go to the <span class="gui">Applications</span> tab and
 check that your application is not muted.</p>
</div></div>
</div></div>
<div id="speakers" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Check that the speakers are turned on and connected properly</span></h2></div>
<div class="region"><div class="contents">
<p class="p">If your computer has external speakers, make sure that they are turned on
 and that the volume is turned up. Make sure that the speaker cable is securely
 plugged into the "output" audio socket on the back of the computer. This socket
 is usually light green in color.</p>
<p class="p">Some sound cards are able to switch which socket they use for output (to the
 speakers) and input (from a microphone, for instance). The output socket may be
 different when running Linux than on Windows or Mac OS. Try connecting the
 speaker cable to the different audio sockets on the computer in turn to see if
 that works.</p>
<p class="p">A final thing to check is that the audio cable is securely plugged into the
 back of the speakers. Some speakers have more than one input too.</p>
</div></div>
</div></div>
<div id="device" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Check that the right sound device is selected</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Some computers have multiple "sound devices" installed. Some of these are
 capable of outputting sound and some are not, so you should check that you have
 the correct one selected. This might involve some trial-and-error to choose the
 right one.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Click the <span class="gui">sound menu</span> in the <span class="gui">menu bar</span> and click <span class="gui">Sound Settings</span>.</p></li>
<li class="steps"><p class="p">In the <span class="gui">Sound</span> window that appears, try selecting a different output from the <span class="gui">Play sound through</span> list.</p></li>
<li class="steps"><p class="p">For the selected device, click <span class="gui">Test Sound</span>.  In the pop-up window, click the
  button for each speaker. Each button will speak its position only to the channel
  corresponding to that speaker.</p></li>
<li class="steps"><p class="p">If that doesn't work, you might want to try doing the same for any other
 devices that are listed.</p></li>
</ol></div></div></div>
</div></div>
</div></div>
<div id="hardware-detected" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Check that the sound card was detected properly</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Your sound card may not have been detected properly. If this has happened,
 your computer will think that it isn't able to play sound. A possible reason
 for the card not being detected properly is that the drivers for the card are
 not installed.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Go to the <span class="link"><a href="unity-dash-intro.html" title="Hitta program, filer, musik och annat med Dash">Dash</a></span> and open the Terminal.</p></li>
<li class="steps"><p class="p">Type <span class="cmd">aplay -l</span> and press <span class="key"><kbd>Enter</kbd></span>.</p></li>
<li class="steps"><p class="p">A list of devices will be shown. If there are no <span class="gui">playback hardware
 devices</span>, your sound card has not been detected.</p></li>
</ol></div></div></div>
<p class="p">If your sound card is not detected, you may need to manually install the
 drivers for it. How you do this will depend on the card you have.</p>
<p class="p">You can see what sound card you have by using the <span class="cmd">lspci</span> command
 in the <span class="app">Terminal</span>. You can get more complete results if you run <span class="cmd">lspci</span> as
 <span class="link"><a href="user-admin-explain.html" title="How do administrative privileges work?">superuser</a></span>; enter <span class="cmd">sudo lspci</span>
 and type your password. See if an
 <span class="em">audio controller</span> or <span class="em">audio device</span> is listed—it should have the
 sound card's make and model number. <span class="cmd">sudo lspci -v</span> will show a list with
 more detailed information.</p>
<p class="p">You may be able to find and install drivers for your card by searching the Internet. Otherwise, you can <span class="link"><a href="report-ubuntu-bug.html" title="Rapportera ett problem i Ubuntu">file a bug</a></span>.</p>
<p class="p">If you can't get drivers for your sound card, you might prefer to buy a new
 sound card. You can get sound cards that can be installed inside the computer
 and external USB sound cards.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="sound-broken.html" title="Sound problems">Sound problems</a><span class="desc"> — Troubleshoot problems like having no sound or having poor sound quality.</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
