<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Användarkonton</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Användarkonton</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Varje person som använder datorn bör ha ett eget användarkonto. Detta låter dem ha sina filer åtskilda från dina samt att ha egna inställningar. Det är också mer säkert. Du kan bara komma åt ett annat användarkonto om du känner till lösenordet.</p></div>
<div id="manage" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Hantera användarkonton</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-add.html" title="Lägg till ett nytt användarkonto"><span class="title">Lägg till ett nytt användarkonto</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till nya användare så att andra personer kan logga in på datorn.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="shell-guest-session.html" title="Starta en begränsad gästsession"><span class="title">Starta en begränsad gästsession</span><span class="linkdiv-dash"> — </span><span class="desc">Låt en vän eller kollega låna din dator på ett säkert sätt.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-delete.html" title="Ta bort ett användarkonto"><span class="title">Ta bort ett användarkonto</span><span class="linkdiv-dash"> — </span><span class="desc">Ta bort användare som inte längre använder din dator.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-changepicture.html" title="Ändra ditt foto på inloggningsskärmen"><span class="title">Ändra ditt foto på inloggningsskärmen</span><span class="linkdiv-dash"> — </span><span class="desc">Lägg till din bild på inloggnings- och användarskärmarna.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="passwords" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Lösenord</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-forgottenpassword.html" title="Jag har glömt mitt lösenord!"><span class="title">Jag har glömt mitt lösenord!</span><span class="linkdiv-dash"> — </span><span class="desc">Avancerade tekniker för att återställa ditt lösenord.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-changepassword.html" title="Välj ditt lösenord"><span class="title">Välj ditt lösenord</span><span class="linkdiv-dash"> — </span><span class="desc">Skydda ditt konto genom att byta lösenord ofta, i dina kontoinställningar.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="user-goodpassword.html" title="Välj ett säkert lösenord"><span class="title">Välj ett säkert lösenord</span><span class="linkdiv-dash"> — </span><span class="desc">Använd längre och mer komplicerade lösenord.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="privileges" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Användarbehörigheter</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="user-admin-explain.html" title="Hur fungerar administratörsbehörighet?"><span class="title">Hur fungerar administratörsbehörighet?</span><span class="linkdiv-dash"> — </span><span class="desc">Du behöver administratörsbehörighet för att ändra viktiga delar i ditt system.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="user-admin-problems.html" title="Problem som orsakas av administratörsbegränsningar"><span class="title">Problem som orsakas av administratörsbegränsningar</span><span class="linkdiv-dash"> — </span><span class="desc">Du kan bara göra vissa saker, som att installera program, om du har administratörsbehörighet.</span></a></div>
</div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="user-admin-change.html" title="Ändra vem som har administratörsbehörighet"><span class="title">Ändra vem som har administratörsbehörighet</span><span class="linkdiv-dash"> — </span><span class="desc">Du kan ändra vilka användare som tillåts göra ändringar för systemet genom att ge dem administratörsbehörighet.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html" title="Mus">mus</a></span>, <span class="link"><a href="prefs-display.html" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html" title="Användarkonton">användarkonton</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
