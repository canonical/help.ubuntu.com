<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Sortera filer och mappar</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="files.html" title="Filer, mappar och sökning">Filer</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Sortera filer och mappar</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan sortera filer på olika sätt i en mapp, till exempel genom att sortera dem efter datum eller filstorlek. Se <span class="link"><a href="#ways" title="Olika sätt att sortera filer">Olika sätt att sortera filer</a></span> nedan för en lista över vanliga sätt att sortera filer. Se <span class="link"><a href="nautilus-views.html" title="Visningsinställningar i Filer">Visningsinställningar i <span class="app">Filer</span></a></span> för information om hur du ändrar standardsorteringen.</p>
<p class="p">Sättet du sorterar filer beror på <span class="em">mappvyn</span> som du använder. Du kan ändra den aktuella vyn via list- eller ikonknapparna i verktygsfältet.</p>
</div>
<div id="icon-view" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Ikonvy</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att sortera filer på ett annat sätt, klicka på <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="nedåtknappen"></span></span>i verktygsfältet och välj <span class="gui">Efter namn</span>, <span class="gui">Efter storlek</span>, <span class="gui">Efter typ</span> eller <span class="gui">Efter ändringsdatum</span>.</p>
<p class="p">Som ett exempel, om du väljer <span class="gui">Efter namn</span> kommer filerna att sorteras efter deras namn i alfabetisk ordning. Se <span class="link"><a href="#ways" title="Olika sätt att sortera filer">Olika sätt att sortera filer</a></span> för ytterligare alternativ.</p>
<p class="p">Du kan sortera i omvänd ordning genom att välja <span class="gui">Omvänd ordning</span> från den utfällbara menyn.</p>
</div></div>
</div></div>
<div id="list-view" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Listvy</span></h2></div>
<div class="region"><div class="contents">
<p class="p">För att sortera filer i en annan ordning, klicka på en av kolumnrubrikerna i filhanteraren. Till exempel, klicka på <span class="gui">Typ</span> för att sortera efter filtyp. Klicka på kolumnrubriken igen för att sortera i omvänd ordning.</p>
<p class="p">I listvyn kan du visa kolumner med fler attribut och sortera efter dessa kolumner. Klicka på <span class="media"><span class="media media-image"><img src="figures/go-down.png" class="media media-inline" alt="nedåtknappen"></span></span> i verktygsfältet, välj <span class="gui">Synliga kolumner</span> och välj vilka kolumner du vill ska vara synliga. Du kommer sedan kunna sortera efter dessa kolumner. Se <span class="link"><a href="nautilus-list.html" title="Inställningar för filhanterarens listkolumner">Inställningar för filhanterarens listkolumner</a></span> för beskrivningar av tillgängliga kolumner.</p>
</div></div>
</div></div>
<div id="ways" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Olika sätt att sortera filer</span></h2></div>
<div class="region"><div class="contents"><div class="terms"><div class="inner"><div class="region"><dl class="terms">
<dt class="terms">Efter namn</dt>
<dd class="terms"><p class="p">Sorterar alfabetiskt efter namnet på filen.</p></dd>
<dt class="terms">Efter storlek</dt>
<dd class="terms"><p class="p">Sorterar efter filens storlek (hur mycket diskutrymme den tar upp). Sorterar från minsta till största som standard.</p></dd>
<dt class="terms">Efter typ</dt>
<dd class="terms"><p class="p">Sorterar alfabetiskt efter filtyp. Filer av samma typ grupperas tillsammans, och sorteras sedan efter namn.</p></dd>
<dt class="terms">Efter ändringsdatum</dt>
<dd class="terms"><p class="p">Sorterar efter tid och datum när en fil senast ändrades. Sorterar som standard från äldst till nyast.</p></dd>
</dl></div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="files.html" title="Filer, mappar och sökning">Filer, mappar och sökning</a><span class="desc"> — <span class="link"><a href="files-search.html" title="Sök efter filer">Sök</a></span>, <span class="link"><a href="files-delete.html" title="Ta bort filer och mappar">radera filer</a></span>, <span class="link"><a href="files.html#backup" title="Säkerhetskopiering">säkerhetskopior</a></span>, <span class="link"><a href="files.html#removable" title="Flyttbara enheter och externa diskar">externa diskar</a></span>, <span class="link"><a href="files.html#documents" title="Dokument">dokument</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
