<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>iSCSI Initiator</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = "index.html.en";
        } else {
                window.location = href.replace(/\.html.*/, ".html.en");
        }
         return false;
      }
      function browserPreferredLanguage() {
        var href = window.location.href;
        if (href.slice(-1) == "/") {
                window.location = href;
        } else {
                window.location = href.replace(/\.html.*/, ".html");
        }
        return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../18.04" class="trail">Ubuntu 18.04</a> » <a class="trail" href="index.html.sv" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="file-servers.html.sv" title="Filservrar">Filservrar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="network-file-system.html.sv" title="Nätverksfilsystem (NFS)">Föregående</a><a class="nextlinks-next" href="cups.html.sv" title="CUPS - Skrivarserver">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">iSCSI Initiator</h1></div>
<div class="region">
<div class="contents">
<p class="para">
      <span class="em emphasis">iSCSI</span> (Internet Small Computer System Interface) is a protocol that allows SCSI commands to be transmitted over a network.
      Typically iSCSI is implemented in a SAN (Storage Area Network) to allow servers to access a large store of hard drive space.  The iSCSI protocol
      refers to clients as <span class="em emphasis">initiators</span> and iSCSI servers as <span class="em emphasis">targets</span>.
      </p>
<p class="para">
      Ubuntu Server can be configured as both an iSCSI initiator and a target.  This guide provides commands and configuration options to setup an iSCSI
      initiator.  It is assumed that you already have an iSCSI target on your local network and have the appropriate rights to connect to it.  The 
      instructions for setting up a target vary greatly between hardware providers, so consult your vendor documentation to configure your specific 
      iSCSI target.
      </p>
</div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="iscsi-initiator.html.sv#iscsi-initiator-install" title="iSCSI Initiator Install">iSCSI Initiator Install</a></li>
<li class="links"><a class="xref" href="iscsi-initiator.html.sv#iscsi-initiator-config" title="iSCSI Initiator Configuration">iSCSI Initiator Configuration</a></li>
<li class="links"><a class="xref" href="iscsi-initiator.html.sv#iscsi-initiator-references" title="Referenser">Referenser</a></li>
</ul></div>
<div class="sect2 sect" id="iscsi-initiator-install"><div class="inner">
<div class="hgroup"><h2 class="title">iSCSI Initiator Install</h2></div>
<div class="region"><div class="contents">
<p class="para">
        To configure Ubuntu Server as an iSCSI initiator install the <span class="app application">open-iscsi</span> package.  In a terminal enter:
        </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo apt install open-iscsi</span>
</pre></div>
</div></div>
</div></div>
<div class="sect2 sect" id="iscsi-initiator-config"><div class="inner">
<div class="hgroup"><h2 class="title">iSCSI Initiator Configuration</h2></div>
<div class="region"><div class="contents">
<p class="para">
        Once the <span class="app application">open-iscsi</span> package is installed, edit <span class="file filename">/etc/iscsi/iscsid.conf</span> changing the following:
        </p>
<div class="code"><pre class="contents ">node.startup = automatic
</pre></div>
<p class="para">
        You can check which targets are available by using the <span class="app application">iscsiadm</span> utility.  Enter the following in a terminal:
        </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo iscsiadm -m discovery -t st -p 192.168.0.10</span>
</pre></div>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist"><p class="para"><span class="em emphasis">-m:</span> determines the mode that iscsiadm executes in.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">-t:</span> specifies the type of discovery.</p></li>
<li class="list itemizedlist"><p class="para"><span class="em emphasis">-p:</span> option indicates the target IP address.</p></li>
</ul></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
          <p class="para">
          Change example <span class="em emphasis">192.168.0.10</span> to the target IP address on your network.
          </p>
        </div></div></div></div>
<p class="para">
        If the target is available you should see output similar to the following:
        </p>
<div class="screen"><pre class="contents "><span class="output computeroutput">
192.168.0.10:3260,1 iqn.1992-05.com.emc:sl7b92030000520000-2
</span>
</pre></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
          <p class="para">
          The <span class="em emphasis">iqn</span> number and IP address above will vary depending on your hardware.
          </p>
        </div></div></div></div>
<p class="para">
        You should now be able to connect to the iSCSI target, and depending on your target 
        setup you may have to enter user credentials.  Login to the iSCSI node: 
        </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo iscsiadm -m node --login</span>
</pre></div>
<p class="para">
        Check to make sure that the new disk has been detected using <span class="app application">dmesg</span>:
        </p>
<div class="screen"><pre class="contents "><span class="cmd command">dmesg | grep sd</span>
<span class="output computeroutput">
[    4.322384] sd 2:0:0:0: Attached scsi generic sg1 type 0
[    4.322797] sd 2:0:0:0: [sda] 41943040 512-byte logical blocks: (21.4 GB/20.0 GiB)
[    4.322843] sd 2:0:0:0: [sda] Write Protect is off
[    4.322846] sd 2:0:0:0: [sda] Mode Sense: 03 00 00 00
[    4.322896] sd 2:0:0:0: [sda] Cache data unavailable
[    4.322899] sd 2:0:0:0: [sda] Assuming drive cache: write through
[    4.323230] sd 2:0:0:0: [sda] Cache data unavailable
[    4.323233] sd 2:0:0:0: [sda] Assuming drive cache: write through
[    4.325312]  sda: sda1 sda2 &lt; sda5 &gt;
[    4.325729] sd 2:0:0:0: [sda] Cache data unavailable
[    4.325732] sd 2:0:0:0: [sda] Assuming drive cache: write through
[    4.325735] sd 2:0:0:0: [sda] Attached SCSI disk
[ 2486.941805] sd 4:0:0:3: Attached scsi generic sg3 type 0
[ 2486.952093] sd 4:0:0:3: [sdb] 1126400000 512-byte logical blocks: (576 GB/537 GiB)
[ 2486.954195] sd 4:0:0:3: [sdb] Write Protect is off
[ 2486.954200] sd 4:0:0:3: [sdb] Mode Sense: 8f 00 00 08
[ 2486.954692] sd 4:0:0:3: [sdb] Write cache: disabled, read cache: enabled, doesn't
 support DPO or FUA
[ 2486.960577]  sdb: sdb1
[ 2486.964862] sd 4:0:0:3: [sdb] Attached SCSI disk
</span>
</pre></div>
<p class="para">
        In the output above <span class="em emphasis">sdb</span> is the new iSCSI disk.  Remember this is just an example; 
        the output you see on your screen will vary.
        </p>
<p class="para">
        Next, create a partition, format the file system, and mount the new iSCSI disk.  In a terminal enter:
        </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo fdisk /dev/sdb</span>
<span class="cmd command">n</span>
<span class="cmd command">p</span>
<span class="cmd command">enter</span>
<span class="cmd command">w</span>
</pre></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents">
          <p class="para">
          The above commands are from inside the <span class="app application">fdisk</span> utility; see <span class="cmd command">man fdisk</span> 
          for more detailed instructions.  Also, the <span class="app application">cfdisk</span> utility is sometimes more user friendly.
          </p>
        </div></div></div></div>
<p class="para">
        Now format the file system and mount it to <span class="file filename">/srv</span> as an example:
        </p>
<div class="screen"><pre class="contents "><span class="cmd command">sudo mkfs.ext4 /dev/sdb1</span>
<span class="cmd command">sudo mount /dev/sdb1 /srv</span>
</pre></div>
<p class="para">
        Finally, add an entry to <span class="file filename">/etc/fstab</span> to mount the iSCSI drive during boot:
        </p>
<div class="code"><pre class="contents ">/dev/sdb1       /srv        ext4    defaults,auto,_netdev 0 0
</pre></div>
<p class="para">
        It is a good idea to make sure everything is working as expected by rebooting the server.
        </p>
</div></div>
</div></div>
<div class="sect2 sect" id="iscsi-initiator-references"><div class="inner">
<div class="hgroup"><h2 class="title">Referenser</h2></div>
<div class="region"><div class="contents">
<p class="para">
        <a href="http://www.open-iscsi.com/" class="ulink" title="http://www.open-iscsi.com/">Open-iSCSI Website</a>
        </p>
<p class="para">
        <a href="http://wiki.debian.org/SAN/iSCSI/open-iscsi" class="ulink" title="http://wiki.debian.org/SAN/iSCSI/open-iscsi">Debian Open-iSCSI page</a>
        </p>
</div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="network-file-system.html.sv" title="Nätverksfilsystem (NFS)">Föregående</a><a class="nextlinks-next" href="cups.html.sv" title="CUPS - Skrivarserver">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address
          so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>
          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p>
</div>
</div>
</body>
</html>
