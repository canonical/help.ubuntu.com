<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Klicka, dra eller rulla med styrplattan</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html.sv" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 22.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html.sv" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Klicka, dra eller rulla med styrplattan</span></h1></div>
<div class="region">
<div class="contents pagewide">
<p class="p">Du kan klicka dubbelklicka, dra och rulla genom att enbart använda din styrplatta, utan andra hårdvaruknappar.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p"><span class="link"><a href="touchscreen-gestures.html.sv" title="Använd gester på styrplattor och pekskärmar">Styrplattegester</a></span> diskuteras separat.</p></div></div></div>
</div>
</div>
<section id="tap"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Knacka för att klicka</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="media media-image floatend"><div class="inner"><img src="figures/touch-tap.svg" class="media media-block" alt=""></div></div>
<p class="p">Du kan knacka på din styrplatta för att klicka istället för att använda en knapp.</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">För att klicka, tryck på styrplattan.</p></li>
<li class="list"><p class="p">För att dubbelklicka, tryck två gånger.</p></li>
<li class="list"><p class="p">För att dra ett objekt, dubbeltryck; men lyft inte fingret efteråt. Dra objektet dit du vill ha det, och lyft sedan fingret för att släppa.</p></li>
<li class="list"><p class="p">Om din styrplatta har stöd för flerfingersknackningar, högerklicka genom att knacka med två fingrar samtidigt. Annars måste du fortfarande använda hårdvaruknapparna för att högerklicka. Se <span class="link"><a href="a11y-right-click.html.sv" title="Simulera ett högerklick">Simulera ett högerklick</a></span> för ett sätt att högerklicka utan en andra musknapp.</p></li>
<li class="list"><p class="p">Om din styrplatta har stöd för flerfingersknackningar, <span class="link"><a href="mouse-middleclick.html.sv" title="Mittenklick">mittenklicka</a></span> genom att knacka med tre fingrar samtidigt.</p></li>
</ul></div></div></div>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">När du trycker eller drar med flera fingrar, se till att dina fingrar är tillräckligt långt från varandra. Om dina fingrar hamnar för tätt ihop kan datorn tro att du bara använder ett finger.</p></div></div></div>
</div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">Aktivera Knacka för att klicka</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Mus &amp; styrplatta</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Mus &amp; styrplatta</span> för att öppna panelen.</p></li>
<li class="steps">
<p class="p">I avsnittet <span class="gui">Styrplatta</span>, säkerställ att <span class="gui">Styrplatta</span> är påslaget.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Avsnittet <span class="gui">Styrplatta</span> visas bara om ditt system har en styrplatta.</p></div></div></div>
</div>
</li>
<li class="steps"><p class="p">Slå på <span class="gui">Knacka för att klicka</span>.</p></li>
</ol></div>
</div></div>
</div></div>
</div></section><section id="twofingerscroll"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Tvåfingersrullning</span></h2></div>
<div class="region"><div class="contents pagewide">
<div class="media media-image floatend"><div class="inner"><img src="figures/touch-scroll.svg" class="media media-block" alt=""></div></div>
<p class="p">Du kan rulla via din styrplatta genom att använda två fingrar.</p>
<p class="p">När detta är valt, kommer att knacka och dra med ett finger att fungera som vanligt men om du drar med två fingrar över någon del av styrplattan kommer den att rulla istället. Flytta fingrarna mellan toppen och botten av styrplattan för att rulla upp och ner, eller flytta fingrarna tvärs över styrplattan för att rulla sidledes. Sprid ut dina fingrar. Om dina fingrar är för nära varandra kommer de att se ut som en stor finger för din styrplatta.</p>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Tvåfingersrullning kanske inte fungerar på alla styrplattor.</p></div></div></div>
</div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">Aktivera Tvåfingersrullning</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Mus &amp; styrplatta</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Mus &amp; styrplatta</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">I avsnittet <span class="gui">Styrplatta</span>, säkerställ att <span class="gui">Styrplatta</span> är påslaget.</p></li>
<li class="steps"><p class="p">Slå på <span class="gui">Tvåfingersrullning</span>.</p></li>
</ol></div>
</div></div>
</div></div>
</div></section><section id="contentsticks"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Naturlig rullning</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Du kan dra innehåll som om du flyttade en fysisk bit papper via styrplattan.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html.sv#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Mus &amp; styrplatta</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Mus &amp; styrplatta</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">I avsnittet <span class="gui">Styrplatta</span>, säkerställ att <span class="gui">Styrplatta</span> är påslaget.</p></li>
<li class="steps"><p class="p">Slå på <span class="gui">Naturlig rullning</span>.</p></li>
</ol></div></div></div>
<div class="note" title="Anteckning">
<svg width="24" height="24" version="1.1">
 <path class="yelp-svg-fill" d="m4 3h16c0.554 0 1 0.446 1 1v11h-6v6h-11c-0.554 0-1-0.446-1-1v-16c0-0.554 0.446-1 1-1z"></path>
 <path class="yelp-svg-fill" d="m17 16h4l-5 5v-4c0-0.554 0.446-1 1-1z"></path>
</svg><div class="inner"><div class="region"><div class="contents"><p class="p">Denna funktion kallas också <span class="em">Omvänd rullning</span>.</p></div></div></div>
</div>
</div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="mouse.html.sv" title="Mus, styrplatta &amp; pekskärm">Mus, styrplatta &amp; pekskärm</a><span class="desc"> — Justera beteendet hos pekdon så att de uppfyller dina personliga krav.</span>
</li></ul></div>
</div></div></div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
