<?xml version="1.0" encoding="utf-8"?>
<ns0:svg xmlns:dc="http://purl.org/dc/elements/1.1/" xmlns:ns0="http://www.w3.org/2000/svg" xmlns:ns1="http://www.inkscape.org/namespaces/inkscape" xmlns:ns2="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd" xmlns:ns3="http://www.openswatchbook.org/uri/2009/osb" xmlns:ns4="http://www.w3.org/1999/xlink" xmlns:ns6="http://creativecommons.org/ns#" xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#" height="500" id="svg10075" version="1.1" width="840" ns2:docname="gs-go-online2.svg" ns1:version="0.92.4 5da689c313, 2019-01-14">
  <ns0:defs id="defs10077">
    <ns0:linearGradient id="linearGradient14901" ns1:collect="always">
      <ns0:stop id="stop14903" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop14905" offset="1" style="stop-color:#000000;stop-opacity:0;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="RHEL7" ns3:paint="gradient">
      <ns0:stop id="stop13323" offset="0" style="stop-color:#a3dbe8;stop-opacity:1;"/>
      <ns0:stop id="stop13325" offset="1" style="stop-color:#a3dbe8;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="GNOME" ns3:paint="gradient">
      <ns0:stop id="stop11074" offset="0" style="stop-color:#eeedec;stop-opacity:1;"/>
      <ns0:stop id="stop11076" offset="1" style="stop-color:#eeedec;stop-opacity:1"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="BLANK" ns3:paint="gradient">
      <ns0:stop id="stop7012" offset="0" style="stop-color:#eeedec;stop-opacity:0;"/>
      <ns0:stop id="stop7014" offset="1" style="stop-color:#eeedec;stop-opacity:0"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(1.1834379,0,0,0.896461,5.7016703,415.60382)" gradientUnits="userSpaceOnUse" id="linearGradient7064" x1="-18.33782" x2="713.42853" y1="490.54935" y2="490.54935" ns1:collect="always" ns4:href="#GNOME"/>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient5885" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient5716">
      <ns0:stop id="stop5718" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient17441" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716"/>
    <ns0:linearGradient id="linearGradient17443">
      <ns0:stop id="stop17445" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop17447" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient3962-1-1-9-5-4-2">
      <ns0:stop id="stop3964-5-0-1-9-6-6" offset="0.0000000" style="stop-color: rgb(211, 233, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4134-0-8-0-8-6-6" offset="0.15517241" style="stop-color: rgb(243, 249, 255); stop-opacity: 1;"/>
      <ns0:stop id="stop4346-9-1-1-2-3-4" offset="0.63108921" style="stop-color: rgb(55, 100, 151); stop-opacity: 1;"/>
      <ns0:stop id="stop6610-2-9-0-2-7" offset="0.81554461" style="stop-color: rgb(39, 62, 93); stop-opacity: 1;"/>
      <ns0:stop id="stop3966-7-2-7-7-1-3" offset="1" style="stop-color: rgb(82, 110, 165); stop-opacity: 1;"/>
    </ns0:linearGradient>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68893" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:linearGradient id="linearGradient6868-5-7-5-4-3" ns1:collect="always">
      <ns0:stop id="stop6870-84-7-0-1-8" offset="0" style="stop-color: rgb(0, 0, 0); stop-opacity: 1;"/>
      <ns0:stop id="stop6872-0-5-0-7-1" offset="1" style="stop-color: rgb(0, 0, 0); stop-opacity: 0;"/>
    </ns0:linearGradient>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68891" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68897" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68895" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68901" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68899" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68905" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68903" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68909" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68907" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68913" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68911" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68917" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68915" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68921" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68919" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68925" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:radialGradient cx="24.881451" cy="22.999987" fx="24.881451" fy="22.999987" gradientTransform="matrix(1,0,0,0.931606,0,1.57305)" gradientUnits="userSpaceOnUse" id="radialGradient68923" r="19.18985" ns1:collect="always" ns4:href="#linearGradient6868-5-7-5-4-3"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath56767">
      <ns0:path d="m 228.45991,29.202459 833.57379,0 0,290.286071 c -330.23641,0 -408.68316,175.76954 -833.57379,175.76954 z" id="path56769" style="color:#000000;fill:#babdb6;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:nodetypes="ccccc" ns1:connector-curvature="0"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath14882">
      <ns0:path d="m 2728,390 a 482,482 0 1 1 -964,0 482,482 0 1 1 964,0 z" id="path14884" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:8.72566223;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(0.35527386,0,0,0.35527386,119.03054,9.4159878)" ns2:cx="2246" ns2:cy="390" ns2:rx="482" ns2:ry="482" ns2:type="arc"/>
    </ns0:clipPath>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient14907" x1="532.43353" x2="532.43353" y1="187.53497" y2="314.62036" ns1:collect="always" ns4:href="#linearGradient14901"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9">
      <ns0:rect height="6.3750005" id="rect6281-1-9" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4">
      <ns0:rect height="5.21591" id="rect6267-1-9" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81">
      <ns0:rect height="4.8734746" id="rect6261-6-6" style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-2-7-1">
      <ns0:rect height="6.3750005" id="rect6281-3-4-6-6" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-1-4-3">
      <ns0:rect height="5.21591" id="rect6267-6-9-5-5" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-3-9">
      <ns0:rect height="4.8734746" id="rect6261-4-5-4" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25942">
      <ns0:rect height="6.3750005" id="rect25944" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25946">
      <ns0:rect height="5.21591" id="rect25948" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25950">
      <ns0:rect height="4.8734746" id="rect25952" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-9-6-0">
      <ns0:rect height="6.3750005" id="rect6281-3-1-6-2" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-6-4-2-8">
      <ns0:rect height="5.21591" id="rect6267-6-9-19-7-4" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-8-2-8-7-5">
      <ns0:rect height="4.8734746" id="rect6261-4-9-2-7-6-1" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25960">
      <ns0:rect height="6.3750005" id="rect25962" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25964">
      <ns0:rect height="5.21591" id="rect25966" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25968">
      <ns0:rect height="4.8734746" id="rect25970" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25972">
      <ns0:rect height="6.3750005" id="rect25974" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25976">
      <ns0:rect height="5.21591" id="rect25978" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25980">
      <ns0:rect height="4.8734746" id="rect25982" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25984">
      <ns0:rect height="6.3750005" id="rect25986" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25988">
      <ns0:rect height="5.21591" id="rect25990" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25992">
      <ns0:rect height="4.8734746" id="rect25994" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath25996">
      <ns0:rect height="6.3750005" id="rect25998" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath26000">
      <ns0:rect height="5.21591" id="rect26002" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath26004">
      <ns0:rect height="4.8734746" id="rect26006" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath24971-0">
      <ns0:rect height="93" id="rect24973-5" style="color:#000000;fill:none;stroke:#000000;stroke-width:2;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="276" x="624" y="-354.29291"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-2-7">
      <ns0:rect height="6.3750005" id="rect6281-3-4-6" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-1-4">
      <ns0:rect height="5.21591" id="rect6267-6-9-5" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-3">
      <ns0:rect height="4.8734746" id="rect6261-4-5" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:mask id="mask12112-0-6-5-3-8-1-7" maskUnits="userSpaceOnUse">
      <ns0:rect height="16" id="rect12114-2-9-0-8-2-5-6" style="fill:url(#radialGradient12116-6-2-9-3-0-9-9);fill-opacity:1;stroke:none" width="221" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient cx="128.5" cy="442" fx="128.5" fy="442" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" gradientUnits="userSpaceOnUse" id="radialGradient12116-6-2-9-3-0-9-9" r="110.5" ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-5-5"/>
    <ns0:linearGradient id="linearGradient12104-5-1-5-6-8-5-5" ns1:collect="always">
      <ns0:stop id="stop12106-3-0-0-5-2-4-1" offset="0" style="stop-color:#cccccc;stop-opacity:1;"/>
      <ns0:stop id="stop12108-4-0-4-9-5-8-15" offset="1" style="stop-color:#cccccc;stop-opacity:0;"/>
    </ns0:linearGradient>
    <ns0:clipPath id="clipPath4201-6-8-5-59">
      <ns0:path d="m 101,177 0,5 2,0 0,2 1,0 0,-4 7,0 0,4 1,0 0,-2 2,0 0,-5 -13,0 z" id="path4203-1-2-5-0" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns1:connector-curvature="0"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6279-6-9-6">
      <ns0:rect height="6.3750005" id="rect6281-3-1-6" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6265-33-6-4-2">
      <ns0:rect height="5.21591" id="rect6267-6-9-19-7" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath id="clipPath6259-6-8-2-8-7">
      <ns0:rect height="4.8734746" id="rect6261-4-9-2-7-6" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:mask id="mask12112-0-6-5-3-8-3-7" maskUnits="userSpaceOnUse">
      <ns0:rect height="16" id="rect12114-2-9-0-8-2-6-5" style="fill:url(#radialGradient12116-6-2-9-3-0-75-13);fill-opacity:1;stroke:none" width="221" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient cx="128.5" cy="442" fx="128.5" fy="442" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" gradientUnits="userSpaceOnUse" id="radialGradient12116-6-2-9-3-0-75-13" r="110.5" ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-7-2"/>
    <ns0:linearGradient id="linearGradient12104-5-1-5-6-8-7-2" ns1:collect="always">
      <ns0:stop id="stop12106-3-0-0-5-2-8-92" offset="0" style="stop-color:#cccccc;stop-opacity:1;"/>
      <ns0:stop id="stop12108-4-0-4-9-5-04-00" offset="1" style="stop-color:#cccccc;stop-opacity:0;"/>
    </ns0:linearGradient>
    <ns0:mask id="mask12112-0-6-5-3-8-0-0" maskUnits="userSpaceOnUse">
      <ns0:rect height="16" id="rect12114-2-9-0-8-2-3-8" style="fill:url(#radialGradient12116-6-2-9-3-0-7-75);fill-opacity:1;stroke:none" width="221" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient cx="128.5" cy="442" fx="128.5" fy="442" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" gradientUnits="userSpaceOnUse" id="radialGradient12116-6-2-9-3-0-7-75" r="110.5" ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-9-1"/>
    <ns0:linearGradient id="linearGradient12104-5-1-5-6-8-9-1" ns1:collect="always">
      <ns0:stop id="stop12106-3-0-0-5-2-3-4" offset="0" style="stop-color:#cccccc;stop-opacity:1;"/>
      <ns0:stop id="stop12108-4-0-4-9-5-0-50" offset="1" style="stop-color:#cccccc;stop-opacity:0;"/>
    </ns0:linearGradient>
    <ns0:mask id="mask12112-0-6-5-3-8-4" maskUnits="userSpaceOnUse">
      <ns0:rect height="16" id="rect12114-2-9-0-8-2-0" style="fill:url(#radialGradient12116-6-2-9-3-0-3);fill-opacity:1;stroke:none" width="221" x="16.5" y="434"/>
    </ns0:mask>
    <ns0:radialGradient cx="128.5" cy="442" fx="128.5" fy="442" gradientTransform="matrix(1,0,0,0.07239819,-1.5,410)" gradientUnits="userSpaceOnUse" id="radialGradient12116-6-2-9-3-0-3" r="110.5" ns1:collect="always" ns4:href="#linearGradient12104-5-1-5-6-8-77"/>
    <ns0:linearGradient id="linearGradient12104-5-1-5-6-8-77" ns1:collect="always">
      <ns0:stop id="stop12106-3-0-0-5-2-87" offset="0" style="stop-color:#cccccc;stop-opacity:1;"/>
      <ns0:stop id="stop12108-4-0-4-9-5-7" offset="1" style="stop-color:#cccccc;stop-opacity:0;"/>
    </ns0:linearGradient>
    <ns0:linearGradient id="linearGradient14901-1" ns1:collect="always">
      <ns0:stop id="stop14903-7" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop14905-2" offset="1" style="stop-color:#000000;stop-opacity:0;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientTransform="matrix(0.75098334,0,0,0.75098334,-170.84871,-42.430559)" gradientUnits="userSpaceOnUse" id="linearGradient27012" x1="532.43353" x2="532.43353" y1="187.53497" y2="314.62036" ns1:collect="always" ns4:href="#linearGradient14901-1"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-9">
      <ns0:rect height="6.3750005" id="rect6281-1-9-8" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4">
      <ns0:rect height="5.21591" id="rect6267-1-9-6" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2">
      <ns0:rect height="4.8734746" id="rect6261-6-6-7" style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-6-1">
      <ns0:rect height="6.3750005" id="rect6281-3-1" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-33-4">
      <ns0:rect height="5.21591" id="rect6267-6-5" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-6-4">
      <ns0:rect height="4.8734746" id="rect6261-4-9" style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath32041">
      <ns0:rect height="6.3750005" id="rect32043" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath32045">
      <ns0:rect height="5.21591" id="rect32047" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-6-8-25-4">
      <ns0:rect height="4.8734746" id="rect6261-4-9-24-2" style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-6-1-4-5">
      <ns0:rect height="6.3750005" id="rect6281-3-0-3-5" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-33-6-5-1-3">
      <ns0:rect height="5.21591" id="rect6267-6-9-1-4-8" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-6-8-2-1-6-6">
      <ns0:rect height="4.8734746" id="rect6261-4-9-2-0-9-0" style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
    <ns0:filter color-interpolation-filters="sRGB" height="1.1308649" id="filter5601" width="1.2058235" x="-0.10291173" y="-0.065432459" ns1:collect="always">
      <ns0:feGaussianBlur id="feGaussianBlur5603" stdDeviation="0.610872" ns1:collect="always"/>
    </ns0:filter>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient48287" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716-6"/>
    <ns0:linearGradient id="linearGradient5716-6">
      <ns0:stop id="stop5718-7" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop5720-7" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient48289" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716-6"/>
    <ns0:linearGradient id="linearGradient33938">
      <ns0:stop id="stop33940" offset="0" style="stop-color:#000000;stop-opacity:1;"/>
      <ns0:stop id="stop33942" offset="1" style="stop-color:#484848;stop-opacity:1;"/>
    </ns0:linearGradient>
    <ns0:linearGradient gradientUnits="userSpaceOnUse" id="linearGradient33948" x1="29.089951" x2="33.971455" y1="11.772627" y2="9.7093649" ns1:collect="always" ns4:href="#linearGradient5716-6"/>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6279-7-9-7">
      <ns0:rect height="6.3750005" id="rect6281-1-9-2" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="3.8250003" x="26.85" y="220.75"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6265-3-4-4-0">
      <ns0:rect height="5.21591" id="rect6267-1-9-2" style="color:#bebebe;fill:#bebebe;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="2.8977277" x="26.96591" y="221.32954"/>
    </ns0:clipPath>
    <ns0:clipPath clipPathUnits="userSpaceOnUse" id="clipPath6259-8-81-2-5">
      <ns0:rect height="4.8734746" id="rect6261-6-6-2" style="color:#bebebe;fill:#bebebe;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible" width="1.8762827" x="26.998718" y="221.50153"/>
    </ns0:clipPath>
  </ns0:defs>
  <ns2:namedview bordercolor="#666666" borderlayer="true" borderopacity="1.0" fit-margin-bottom="0" fit-margin-left="0" fit-margin-right="0" fit-margin-top="0" height="0px" id="base" pagecolor="#eeeeec" showgrid="false" width="0px" ns1:current-layer="g26899" ns1:cx="0.46369647" ns1:cy="354.43398" ns1:document-units="px" ns1:pageopacity="1" ns1:pageshadow="2" ns1:showpageshadow="false" ns1:window-height="1401" ns1:window-maximized="1" ns1:window-width="2560" ns1:window-x="2560" ns1:window-y="0" ns1:zoom="1">
    <ns1:grid empspacing="5" enabled="true" id="grid17504" snapvisiblegridlinesonly="true" type="xygrid" visible="true"/>
  </ns2:namedview>
  <ns0:metadata id="metadata10080">
    <rdf:RDF>
      <ns6:Work rdf:about="">
        <dc:format>image/svg+xml</dc:format>
        <dc:type rdf:resource="http://purl.org/dc/dcmitype/StillImage"/>
        <dc:title/>
      </ns6:Work>
    </rdf:RDF>
  </ns0:metadata>
  <ns0:g id="layer1" transform="translate(0,-992.3622)" ns2:insensitive="true" ns1:groupmode="layer" ns1:label="bg">
    <ns0:rect height="656" id="background" style="fill:url(#BLANK);" width="866" x="-16" y="855.36218" ns1:label="background"/>
  </ns0:g>
  <ns0:g id="layer2" transform="translate(0,-540)" ns1:groupmode="layer" ns1:label="fg">
    <ns0:g id="g27126" transform="translate(9,-167.29113)">
      <ns0:g id="g15031" transform="translate(-51,24.637831)">
        <ns0:path d="m 137,278 c 0,9.38884 -7.61116,17 -17,17 -9.38884,0 -17,-7.61116 -17,-17 0,-9.38884 7.61116,-17 17,-17 9.38884,0 17,7.61116 17,17 z" id="path15033" style="color:#000000;fill:#000000;fill-opacity:0.27522936;stroke:none;stroke-width:1.06985807;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="translate(2,453.36217)" ns2:cx="120" ns2:cy="278" ns2:rx="17" ns2:ry="17" ns2:type="arc"/>
        <ns0:text id="text15035" style="font-style:normal;font-variant:normal;font-weight:bold;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Bold';text-align:center;letter-spacing:0px;word-spacing:0px;writing-mode:lr-tb;text-anchor:middle;fill:#ffffff;fill-opacity:1;stroke:none" x="122.29289" y="736.36218" xml:space="preserve"><ns0:tspan id="tspan15037" style="font-size:14px;line-height:1.25" x="122.29289" y="736.36218" ns2:role="line">1</ns0:tspan></ns0:text>
      </ns0:g>
      <ns0:g clip-path="none" id="g26899" transform="matrix(0.7432991,0,0,0.7432991,3.7849383,392.29986)">
        <ns0:path d="m 659.42842,512.06341 c -0.7509,0 -1.48468,0.26524 -2.06007,0.84084 l -23.88003,23.88003 -308.21205,0 c -6.5103,0 -11.77184,5.26154 -11.77184,11.77184 l 0,164.46945 427.444,0 0,-164.46945 c 0,-6.5102 -5.2196,-11.77184 -11.7298,-11.77184 l -43.85012,0 -23.88002,-23.88003 c -0.5755,-0.5754 -1.30917,-0.84084 -2.06007,-0.84084 z m -345.92399,348.95104 0,132.47526 c 0,6.51019 5.26154,11.77189 11.77184,11.77189 l 403.94236,0 c 6.5102,0 11.7298,-5.2617 11.7298,-11.77189 l 0,-132.47526 z" id="rect41123-4" style="color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2.93785119;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:nodetypes="sccssccssccscsssscc" ns1:connector-curvature="0"/>
        <ns0:g id="default-pointer-c" style="display:inline" transform="matrix(3.7117385,0,0,3.7117385,441.75165,732.88835)" ns1:label="#g5607">
          <ns0:path d="m 27.135224,2.8483222 0,16.4402338 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 27.135224,2.8483222 z" id="path5567" style="opacity:0.6;color:#000000;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:#000000;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;filter:url(#filter5601);enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
          <ns0:path d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path5565" style="color:#000000;fill:url(#linearGradient48287);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
          <ns0:path d="m 26.604893,2.3179921 0,16.4402329 3.712311,-3.623922 2.12132,4.331029 c 0.519598,1.171377 3.220861,0.229524 2.452777,-1.336875 l -2.099224,-4.496756 4.684582,0 L 26.604893,2.3179921 z" id="path6242" style="color:#000000;fill:url(#linearGradient33948);fill-opacity:1;fill-rule:nonzero;stroke:#ffffff;stroke-width:1;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:10;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:block;overflow:visible;enable-background:accumulate" ns2:nodetypes="cccccccc" ns1:connector-curvature="0"/>
        </ns0:g>
        <ns0:g id="g15062" style="fill:#000000;fill-opacity:1;display:inline" transform="matrix(1.3453534,0,0,1.3453534,332.63788,598.67052)">
          <ns0:g id="g15066" style="fill:#ffffff;fill-opacity:1;display:inline" transform="translate(-81,-317)" ns1:label="status">
            <ns0:g id="g15068" style="fill:#ffffff;fill-opacity:1;display:inline" transform="translate(0,40)">
              <ns0:rect height="2" id="rect15070" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="2.9722719" x="81" y="284"/>
              <ns0:rect height="2" id="rect15072" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="3.0164659" x="93.983536" y="284"/>
            </ns0:g>
            <ns0:g id="g15074" style="fill:#ffffff;fill-opacity:1;display:inline" transform="matrix(0.70710678,-0.70710679,0.70710679,0.70710678,-175.45794,186.40707)">
              <ns0:rect height="2" id="rect15076" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="2.9722719" x="81" y="284"/>
              <ns0:rect height="2" id="rect15078" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="3.0164659" x="93.983536" y="284"/>
            </ns0:g>
            <ns0:g id="g15080" style="fill:#ffffff;fill-opacity:1;display:inline" transform="matrix(0,-1,1,0,-196,414)">
              <ns0:rect height="2" id="rect15082" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="2.9722719" x="81" y="284"/>
              <ns0:rect height="2" id="rect15084" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="3.0164659" x="93.983536" y="284"/>
            </ns0:g>
            <ns0:g id="g15086" style="fill:#ffffff;fill-opacity:1;display:inline" transform="matrix(-0.70710679,-0.70710678,0.70710678,-0.70710679,-49.592928,589.45794)">
              <ns0:rect height="2" id="rect15088" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="2.9722719" x="81" y="284"/>
              <ns0:rect height="2" id="rect15090" rx="0.5625" ry="0.5625" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:new" width="3.0164659" x="93.983536" y="284"/>
            </ns0:g>
            <ns0:path d="m 89.034905,320.9942 c -2.171787,0 -3.946856,1.77507 -3.946856,3.94686 0,2.17178 1.775069,3.97566 3.946856,3.97566 2.171787,0 3.975664,-1.80388 3.975664,-3.97566 0,-2.17179 -1.803877,-3.94686 -3.975664,-3.94686 z m 0,2.01664 c 1.090904,0 1.959023,0.83931 1.959023,1.93022 0,1.0909 -0.868119,1.95902 -1.959023,1.95902 -1.090904,0 -1.930214,-0.86812 -1.930214,-1.95902 0,-1.09091 0.83931,-1.93022 1.930214,-1.93022 z" id="path15092" style="font-size:medium;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;text-indent:0;text-align:start;text-decoration:none;line-height:normal;letter-spacing:normal;word-spacing:normal;text-transform:none;direction:ltr;block-progression:tb;writing-mode:lr-tb;text-anchor:start;baseline-shift:baseline;color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2.16944861;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate;font-family:Sans;-inkscape-font-specification:Sans" ns1:connector-curvature="0"/>
          </ns0:g>
          <ns0:g id="g15094" style="fill:#ffffff;fill-opacity:1" transform="translate(-81,-317)" ns1:label="devices"/>
          <ns0:g id="g15096" style="fill:#ffffff;fill-opacity:1" transform="translate(-81,-317)" ns1:label="apps"/>
          <ns0:g id="g15098" style="fill:#ffffff;fill-opacity:1" transform="translate(-81,-317)" ns1:label="actions"/>
          <ns0:g id="g15100" style="fill:#ffffff;fill-opacity:1" transform="translate(-81,-317)" ns1:label="places"/>
          <ns0:g id="g15102" style="fill:#ffffff;fill-opacity:1" transform="translate(-81,-317)" ns1:label="mimetypes"/>
          <ns0:g id="g15104" style="fill:#ffffff;fill-opacity:1;display:inline" transform="translate(-81,-317)" ns1:label="emblems"/>
          <ns0:g id="g15106" style="fill:#ffffff;fill-opacity:1;display:inline" transform="translate(-81,-317)" ns1:label="categories"/>
        </ns0:g>
        <ns0:rect height="345.7753" id="rect15756" rx="1.8594906" ry="1.7873727" style="color:#000000;fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1.32587242;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(0,1,-1,0,0,0)" width="3.7617662" x="607.55249" y="-720.68964"/>
        <ns0:path d="m 856.7519,116.95945 c 0,2.02705 -1.64325,3.6703 -3.6703,3.6703 -2.02704,0 -3.67029,-1.64325 -3.67029,-3.6703 0,-2.02705 1.64325,-3.6703 3.67029,-3.6703 2.02705,0 3.6703,1.64325 3.6703,3.6703 z" id="path15762" style="fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1;stroke-opacity:1;display:inline" transform="matrix(0,2.6014918,-2.6014918,0,910.14466,-1609.8514)" ns2:cx="853.0816" ns2:cy="116.95945" ns2:rx="3.6702957" ns2:ry="3.6702957" ns2:type="arc"/>
        <ns0:rect height="345.7753" id="rect59830" rx="1.8594906" ry="1.7873727" style="color:#000000;fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1.32587242;stroke-linecap:butt;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(0,1,-1,0,0,0)" width="3.7617662" x="569.88251" y="-720.68964"/>
        <ns0:path d="m 856.7519,116.95945 c 0,2.02705 -1.64325,3.6703 -3.6703,3.6703 -2.02704,0 -3.67029,-1.64325 -3.67029,-3.6703 0,-2.02705 1.64325,-3.6703 3.67029,-3.6703 2.02705,0 3.6703,1.64325 3.6703,3.6703 z" id="path59832" style="fill:#ffffff;fill-opacity:0.99918698;stroke:#000000;stroke-width:1;stroke-opacity:1;display:inline" transform="matrix(0,2.6014918,-2.6014918,0,955.88668,-1647.5213)" ns2:cx="853.0816" ns2:cy="116.95945" ns2:rx="3.6702957" ns2:ry="3.6702957" ns2:type="arc"/>
        <ns0:g id="g5525-4-0" style="fill:#ffffff;fill-opacity:1;display:inline" transform="matrix(1.3453534,0,0,1.3453534,308.37527,269.05896)" ns1:label="audio-speakers">
          <ns0:path d="m 27.433982,218 -3.84375,4.03125 -3.5625,0 0,6.125 3.5625,0 3.9375,3.84375 0.5,-0.0312 0,-13.9375 z" id="path5533-7" style="color:#bebebe;fill:#ffffff;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" ns2:nodetypes="ccccccccc" ns1:connector-curvature="0"/>
          <ns0:path d="m 30.939342,221 2,-2" id="path8311" style="fill:none;stroke:#ffffff;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
          <ns0:path d="m 30.939342,229 2,2" id="path9081" style="fill:none;stroke:#ffffff;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
          <ns0:path d="m 31.939342,225.0202 3.03125,0" id="path9083" style="color:#000000;fill:none;stroke:#ffffff;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;stroke-dashoffset:0;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
          <ns0:rect height="1" id="rect9102" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.0000017" x="29.93936" y="221"/>
          <ns0:rect height="1" id="rect9104" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:2;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="1.0000017" x="29.93936" y="228"/>
        </ns0:g>
        <ns0:rect height="44.396664" id="rect59873" rx="0" ry="0" style="color:#000000;fill:#ffffff;fill-opacity:1;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" width="429.16772" x="312.41132" y="668.62891"/>
        <ns0:text id="text32132" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="366.59216" y="698.00366" xml:space="preserve"><ns0:tspan id="tspan32134" style="font-size:20.56496048px;line-height:1.25" x="366.59216" y="698.00366" ns2:role="line">Trådlöst nätverk</ns0:tspan></ns0:text>
        <ns0:g id="g3944" style="display:inline" transform="matrix(1.3453534,0,0,1.3453534,274.74144,415.70247)" ns1:label="network-wireless-signal-good">
          <ns0:path clip-path="url(#clipPath6279-6-1)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" id="path3743" style="fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" transform="matrix(0,-0.784314,0.784314,0,-128.137,227.059)" ns2:cx="24.9375" ns2:cy="223.9375" ns2:end="7.0685835" ns2:open="true" ns2:rx="3.1875" ns2:ry="3.1875" ns2:start="5.4977871" ns2:type="arc"/>
          <ns0:path clip-path="url(#clipPath6265-33-4)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" id="path3745-5" style="fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" transform="matrix(0,-1.72549,1.72549,0,-338.902,250.529)" ns2:cx="24.9375" ns2:cy="223.9375" ns2:end="7.0685835" ns2:open="true" ns2:rx="3.1875" ns2:ry="3.1875" ns2:start="5.4977871" ns2:type="arc"/>
          <ns0:rect height="16" id="rect3749" style="color:#bebebe;fill:none;stroke:none;stroke-width:1;marker:none;visibility:visible;display:inline;overflow:visible" transform="matrix(0,-1,1,0,0,0)" width="16" x="-212" y="40" ns1:label="audio-volume-high"/>
          <ns0:path d="m 29,209 c 0,0.55228 -0.447715,1 -1,1 -0.552285,0 -1,-0.44772 -1,-1 0,-0.55228 0.447715,-1 1,-1 0.552285,0 1,0.44772 1,1 z" id="path3751" style="fill:#000000;fill-opacity:1;stroke:none;display:inline" transform="matrix(1.5,0,0,1.5,5.5,-105)" ns2:cx="28" ns2:cy="209" ns2:rx="1" ns2:ry="1" ns2:type="arc"/>
          <ns0:path clip-path="url(#clipPath6259-6-8-25-4)" d="m 27.191403,221.6836 c 1.244796,1.24479 1.244796,3.26301 0,4.5078 0,0 0,0 0,0" id="path2937-7" style="opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;display:inline" transform="matrix(0,-2.66667,2.66667,0,-549.666,274)" ns2:cx="24.9375" ns2:cy="223.9375" ns2:end="7.0685835" ns2:open="true" ns2:rx="3.1875" ns2:ry="3.1875" ns2:start="5.4977871" ns2:type="arc"/>
        </ns0:g>
        <ns0:text id="text59875" style="color:#000000;font-style:normal;font-variant:normal;font-weight:normal;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:Cantarell;text-indent:0;text-align:end;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:end;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="698.89441" y="698.00366" xml:space="preserve"><ns0:tspan id="tspan59877" style="font-size:20.56496048px;line-height:1.25" x="698.89441" y="698.00366" ns2:role="line">hemmanätverk</ns0:tspan></ns0:text>
        <ns0:path d="m 726.44385,688.97738 -5.04507,5.04508 -5.04509,-5.04508 z" id="rect12003" style="color:#000000;fill:#000000;fill-opacity:1;stroke:none;stroke-width:3;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" ns2:nodetypes="cccc" ns1:connector-curvature="0"/>
        <ns0:text id="text59897" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="331.61298" y="753.16315" xml:space="preserve"><ns0:tspan id="tspan59899" style="font-size:20.56496048px;line-height:1.25" x="331.61298" y="753.16315" ns2:role="line">Välj nätverk</ns0:tspan></ns0:text>
        <ns0:text id="text59901" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="331.61298" y="796.2146" xml:space="preserve"><ns0:tspan id="tspan59903" style="font-size:20.56496048px;line-height:1.25" x="331.61298" y="796.2146" ns2:role="line">Stäng av</ns0:tspan></ns0:text>
        <ns0:text id="text59905" style="color:#000000;font-style:normal;font-variant:normal;font-weight:500;font-stretch:normal;line-height:0%;font-family:Cantarell;-inkscape-font-specification:'Cantarell Medium';text-indent:0;text-align:start;text-decoration:none;text-decoration-line:none;letter-spacing:normal;word-spacing:normal;text-transform:none;writing-mode:lr-tb;direction:ltr;text-anchor:start;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1px;marker:none;enable-background:accumulate" x="331.61298" y="839.26605" xml:space="preserve"><ns0:tspan id="tspan59907" style="font-size:20.56496048px;line-height:1.25" x="331.61298" y="839.26605" ns2:role="line">Inställningar för trådlösa nätverk</ns0:tspan></ns0:text>
        <ns0:g id="g5525" style="display:inline" transform="matrix(1.3453534,0,0,1.3453534,590.89949,182.95633)" ns1:label="audio-volume-medium">
          <ns0:path d="m 20,222 h 2.484375 L 25.453129,219 26,219.0156 v 11 l -0.475297,8.3e-4 L 22.484375,227 H 20 Z" id="path5533" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:1;marker:none" ns2:nodetypes="ccccccccc" ns1:connector-curvature="0"/>
          <ns0:rect height="16" id="rect5535" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" width="16" x="20" y="217" ns1:label="audio-volume-high"/>
          <ns0:path clip-path="url(#clipPath6279-7-9-7)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" id="path3718-5" style="display:inline;fill:none;stroke:#000000;stroke-width:2.54999995;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" transform="matrix(0.784314,0,0,0.784314,5.94118,48.8628)" ns2:cx="24.9375" ns2:cy="223.9375" ns2:end="0.78539819" ns2:open="true" ns2:rx="3.1875" ns2:ry="3.1875" ns2:start="5.4977871" ns2:type="arc"/>
          <ns0:path clip-path="url(#clipPath6265-3-4-4-0)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" id="path3726-1" style="display:inline;fill:none;stroke:#000000;stroke-width:1.15909004;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" transform="matrix(1.72549,0,0,1.72549,-17.5294,-161.902)" ns2:cx="24.9375" ns2:cy="223.9375" ns2:end="0.78539819" ns2:open="true" ns2:rx="3.1875" ns2:ry="3.1875" ns2:start="5.4977871" ns2:type="arc"/>
          <ns0:path clip-path="url(#clipPath6259-8-81-2-5)" d="m 27.191403,221.6836 a 3.1875,3.1875 0 0 1 0.933597,2.2539 3.1875,3.1875 0 0 1 -0.933597,2.2539" id="path3728-0" style="display:inline;opacity:0.35;fill:none;stroke:#000000;stroke-width:0.75;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" transform="matrix(2.66667,0,0,2.66667,-41,-372.666)" ns2:cx="24.9375" ns2:cy="223.9375" ns2:end="0.78539819" ns2:open="true" ns2:rx="3.1875" ns2:ry="3.1875" ns2:start="5.4977871" ns2:type="arc"/>
        </ns0:g>
        <ns0:g id="g4692-3" style="display:inline" transform="matrix(1.3453534,0,0,1.3453534,591.45102,-450.08783)" ns1:label="system-shutdown">
          <ns0:rect height="16" id="rect10837-3-0" rx="0.14408804" ry="0.15129246" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none;enable-background:new" width="16" x="40" y="688"/>
          <ns0:path d="m 51.52343,689.95141 a 7,7 0 0 1 3.233191,7.87837 7,7 0 0 1 -6.766907,5.17021 7,7 0 0 1 -6.751683,-5.19008 7,7 0 0 1 3.25633,-7.86883" id="path3869-2" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:none;stroke:#000000;stroke-width:2.333606;stroke-linecap:round;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1;marker:none;enable-background:accumulate" transform="matrix(0.85694274,0,0,0.85714276,6.8667487,99.42864)" ns2:cx="48" ns2:cy="696" ns2:end="4.1878597" ns2:open="true" ns2:rx="7" ns2:ry="7" ns2:start="5.239857" ns2:type="arc"/>
          <ns0:path d="m 48,689 v 5" id="path4710" style="fill:none;stroke:#000000;stroke-width:2;stroke-linecap:round;stroke-linejoin:miter;stroke-miterlimit:4;stroke-dasharray:none;stroke-opacity:1" ns2:nodetypes="cc" ns1:connector-curvature="0"/>
        </ns0:g>
        <ns0:path d="m 685.77004,486.8382 -5.04507,5.04509 -5.04508,-5.04509 z" id="rect12003-0" style="color:#000000;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;stroke:none;stroke-width:4.03606033;marker:none;enable-background:accumulate" ns2:nodetypes="cccc" ns1:connector-curvature="0"/>
        <ns0:path d="m 301,405.5 c 0,8.00813 -6.49187,14.5 -14.5,14.5 -8.00813,0 -14.5,-6.49187 -14.5,-14.5 0,-8.00813 6.49187,-14.5 14.5,-14.5 8.00813,0 14.5,6.49187 14.5,14.5 z" id="path59993" style="color:#000000;fill:none;stroke:#ffffff;stroke-width:0.8108108;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(1.6592692,0,0,1.6592692,-113.19122,279.66482)" ns2:cx="286.5" ns2:cy="405.5" ns2:rx="14.5" ns2:ry="14.5" ns2:type="arc"/>
        <ns0:path d="m 301,405.5 c 0,8.00813 -6.49187,14.5 -14.5,14.5 -8.00813,0 -14.5,-6.49187 -14.5,-14.5 0,-8.00813 6.49187,-14.5 14.5,-14.5 8.00813,0 14.5,6.49187 14.5,14.5 z" id="path59995" style="color:#000000;fill:none;stroke:#ffffff;stroke-width:0.8108108;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(1.6592692,0,0,1.6592692,212.38431,279.66482)" ns2:cx="286.5" ns2:cy="405.5" ns2:rx="14.5" ns2:ry="14.5" ns2:type="arc"/>
        <ns0:path d="m 301,405.5 c 0,8.00813 -6.49187,14.5 -14.5,14.5 -8.00813,0 -14.5,-6.49187 -14.5,-14.5 0,-8.00813 6.49187,-14.5 14.5,-14.5 8.00813,0 14.5,6.49187 14.5,14.5 z" id="path59997" style="color:#000000;fill:none;stroke:#ffffff;stroke-width:0.8108108;stroke-miterlimit:4;stroke-opacity:1;stroke-dasharray:none;marker:none;visibility:visible;display:inline;overflow:visible;enable-background:accumulate" transform="matrix(1.6592692,0,0,1.6592692,52.287251,279.66482)" ns2:cx="286.5" ns2:cy="405.5" ns2:rx="14.5" ns2:ry="14.5" ns2:type="arc"/>
        <ns0:g id="g8415" style="display:inline;enable-background:new" transform="matrix(1.3453534,0,0,1.3453534,262.633,236.77047)" ns1:label="network-wired">
          <ns0:rect height="16" id="rect8417" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:none;stroke:none;stroke-width:1;marker:none" width="16" x="241.0002" y="177"/>
          <ns0:rect height="4.9375" id="rect8421" ry="0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate" width="5.0000014" x="241.0002" y="188"/>
          <ns0:rect height="5.0000024" id="rect8425" ry="0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate" width="5.0000014" x="251.0002" y="188"/>
          <ns0:path d="M 2.53125,-8.4687501 V -11.5 H 12.5 v 3.0312499" id="path8427" style="fill:none;stroke:#1e2224;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" transform="translate(241.0002,197)" ns2:nodetypes="cccc" ns1:connector-curvature="0"/>
          <ns0:path d="M 7.5,-11.5 V -15" id="path9198" style="fill:none;stroke:#000000;stroke-width:1px;stroke-linecap:butt;stroke-linejoin:miter;stroke-opacity:1" transform="translate(241.0002,197)" ns1:connector-curvature="0"/>
          <ns0:rect height="5.0000024" id="rect9200" ry="0" style="color:#bebebe;display:inline;overflow:visible;visibility:visible;fill:#000000;fill-opacity:1;fill-rule:nonzero;stroke:none;stroke-width:0;marker:none;enable-background:accumulate" width="5.0000014" x="246.0002" y="178"/>
        </ns0:g>
      </ns0:g>
    </ns0:g>
  </ns0:g>
</ns0:svg>
