�PNG

   IHDR  "   �   �SF�   �zTXtRaw profile type exif  x�mP�� ��?B�q�I�n��k�#%mO���0���:� �e�j���5w�L��Xd� Qzx�C?�R4�[���i����bso��3�^0I}�ʇ8&"w��b�L�6�U��z�B��:�T��XV�޶�;L���9#���0ps��=�Foh�����B���| �-Z9����  �iCCPICC profile  x�}�=H�@�_S�"�q�P����U(B�P+��`r�4iHR\ׂ��Ug]\A����I�EJ�_Rh��q?��{ܽ�F�iV�,�鶙N&�lnU�"�D0Qf�1'I)���{�z�Y���}j�b@@$�e�ioOo��}�(+�*�9�I$~�����ό���<q�X,v����dj�S�1U�)_�z�r��Uj�uO��p^_Y�:�a$��%H���2*��U'�B��>�!�/�K!W��B������w�Var�K
'����B�@��8�ǎ�<������W��'���;����붦��;���!��+i
��~Fߔ"�@��[k�@��J� ��h���}����ۿgZ�� ��r�(˞�  viTXtXML:com.adobe.xmp     <?xpacket begin="﻿" id="W5M0MpCehiHzreSzNTczkc9d"?>
<x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 4.4.0-Exiv2">
 <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
  <rdf:Description rdf:about=""
    xmlns:xmpMM="http://ns.adobe.com/xap/1.0/mm/"
    xmlns:stEvt="http://ns.adobe.com/xap/1.0/sType/ResourceEvent#"
    xmlns:dc="http://purl.org/dc/elements/1.1/"
    xmlns:GIMP="http://www.gimp.org/xmp/"
    xmlns:tiff="http://ns.adobe.com/tiff/1.0/"
    xmlns:xmp="http://ns.adobe.com/xap/1.0/"
   xmpMM:DocumentID="gimp:docid:gimp:c0b80621-8646-41ed-9c2f-f01138adca86"
   xmpMM:InstanceID="xmp.iid:8d85b4d4-a8f6-4d8e-8d6e-bcded0760a92"
   xmpMM:OriginalDocumentID="xmp.did:64c69a6c-a38f-415e-9a2d-7f1e24e3b22e"
   dc:Format="image/png"
   GIMP:API="3.0"
   GIMP:Platform="Linux"
   GIMP:TimeStamp="1679601746723488"
   GIMP:Version="2.99.14"
   tiff:Orientation="1"
   xmp:CreatorTool="GIMP"
   xmp:MetadataDate="2023:03:23T21:02:26+01:00"
   xmp:ModifyDate="2023:03:23T21:02:26+01:00">
   <xmpMM:History>
    <rdf:Seq>
     <rdf:li
      stEvt:action="saved"
      stEvt:changed="/"
      stEvt:instanceID="xmp.iid:54dd0f56-317a-40bf-b548-cdd3f21a30ea"
      stEvt:softwareAgent="GIMP 2.99.14 (Linux)"
      stEvt:when="2023-03-23T21:02:26+01:00"/>
    </rdf:Seq>
   </xmpMM:History>
  </rdf:Description>
 </rdf:RDF>
</x:xmpmeta>
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                                                                                                    
                           
<?xpacket end="w"?>����   	pHYs  �  ��+   tIME�
*==   tEXtComment Created with GIMPW�    IDATx��}w|ŵ�9���_IW�K��.˽a0�M���GB �<�彗BBBIȏ$/�^L5���{o�%K��U���;����^ɶ�Us��~?�ȫݝ��s�̙s0
�Ã=��7_��Dd���
f5��4��9�5������gV �l5��adY� Bi�2���c]���h�-ē|�O�_�� �M����驗��f�t�9	Œ�G,��¿�h2���7���ˊ�Q��A}����V-��O*�}gQ��  6U��E��v��֚���Āx_lp��cg9)��/J����)�x_մ�i缦����Zblܸq��� PU]][S�s>j�Ȣ�"Ɔ�4EDG�=\U cǌ���ADM�<X��P\T<bD�$I'=����]QQ�p88����;V��z��'���g��l�.N�:X\�@���ج��_����Z��}�4Y�l*��ɷIY����}_�!h&3�gӉ�ԩ�<��f?��W�.?��ﶣ ��c�W��{�ZFN/����x���v��m��I]�9��֮:����|�cǎm��h��W^mkk۳g��O<��h۶m���F{{�3�>�w��S�Z��������AD{��}����5k�,_�\Ӵd��k�_T��:XL�?~��+-� ��er�-��6%Ic@O�cE��w��H ��*}��[
�x�Gr�z�"�Ms�cr���u����n�,�_5�-�>���4�V�|i��������?��e,s��7�x �:���j�-,,7=z,����9��������X<6rĈ���斖ښZMӊ��rssu]?t�02�F�cF���;���a���o!b �����(�����_��-�E���Y+���q�-{]��/\���6m��dfe m޲yʔ�K/������g���^�gHL crl p�I}qc 8��S�,?-)=���s��G�~���m�d��]�6*KI\��x�'<�>��
Y^)�ҽ�:!_9����w�'���Q�-!��]T�Zs0z�Q��fg��b���ng��.�u������e��y�NY�zu�ccF�޵k��a9rdݱc�7o��Wo=|�𑚚���+W��w���㣏����3f䈑6�rj���eY����h,VXP @�9�mmm��I�HD�@�֭[�^��eˀ��&N������}釫�&O��t:�6��$�p ��H�iR]�>:Gq�P�;eT���ܔL��ՈrY�kRa������nWw���'�Lc@�q4>�������ѳ晛"ex��Q �m��덶�� �Do>˛� Tkmvƭ�>���qc�*� �p��זm۾����f;A_�\Q���E��E+W���766����s�2erIIIGG�?���ђ�����+�\^\\���n�yy�^����֦(�6��WU"(5J�}��;���0�`iiInn��K���|�g�B�vxoWxF�-�+�����^�-�d<Ԥ�8���T��О�"�:��q (I��ҤT'�W�
�c�V͓~�	4N�� ��XDM�/��Ls�N�zoK��kp�`��;n��+B�8��/�p�K�����+V���-7',�$#bVf��i����\����5Gj|�>�I��D$˲�n/<�Ě��u���r�M���]�p$���,��H��p���|�`�;�;��b�Νx���n���W_[6����/y��-/����������!1����n8�7ʑ�"�Œ��M����,�?{���9��������\�r�8�IOh���M+N�.�^�<߶�&�PPB��=~qS���J���
w�>k���Co��2d@`�9��Ӂ^|�k��:/'��t]���X�n�����c�14/ꪅ���իWO�6���}> 2^�m�DU���z��/]ueQQ!q���LMIٶm{<?t�PQa!",_���o�STT�������/[�hQAA��sϕ$VWW����p�Ǎː�B�d+��$��?�UgX����)�ήp���蒴��z=���Y������/Nu�J��Jֈ��մm��;�m�gi�As���i˶��ݒ"ak�[v�⛫c7���aw*(1p�p�h�U���E�[�^��e9�t��c.���~��ӹs���d���+D����/�`Q�S��C �� �f��������y-�-�m��pr����?���8�͛7o޲e���&L����y��;vt�K.�KKK����p�@$q�\yy�n���s�Y��yy��P���(+++�aC}��`���w�������;�	;^�� v����|[��А��D�9R�ݫ��ƀ��Cq���t �iվ�J�0跅y �#�B1����/����K|k+c�A=?M�=±�>���`T�훱���5�O'TU=XYI�>hAA~JJJSSS�� �4_Ff�d.����EIMM������yyy\����
C�P]}�,�6�-==�a����g�d���u���87PNnNfF��yccc�#���������-8����9ي,�^_�mv[nn���L�����ݯ�}ކ�J�g�9_�ў�v��_��B"��喏D��o�
�'���Mb��c� �Mv�����Q�Nu1������wexXC��j_��}�>��բ��aþF��kꐿ�K��cs!a^��m� হ��t	 :�������N,�aûs1/}ys7[dO�qƶ�l���0��^�4��9�f�?�Y�f,q6ܰ�X�d��K����oݴv�!�y��^:�!�"�0D�e�]�l�����x����3U��-b��z&�b�t<i��	rʯO���[蔻Oy�K+� Nz��Q}��v�o�D�A���훩���t`��TI���I1Y�R�4�>ړN���]ٟ�;	䪍���'$c�q$D" B $f<@D��F��HH@�8p �\�A �Ѥ p��:���x!#�hH]�&GBB�LfM� ���t�o" Ɓ��$�� �� �8 
��$�z� G��+�8p����@"@"4*�u��Dcl/ uan��t D��Oc�ٸ[�N48��#^��Ȉ������8�p�ɑ��F�����Ţ�� �qHt8!'0Ƌ1`�����8 ��	�h�� T�)N%�։�"7�ެ�)4Cc�NDF{��N��˃]�>� ��w" p B��n������iYԻӑ �#$ �eA�$>��#ň$4�Y8PR��Ŧ����qD��1F@$QN�f;p�R4�1[ �`�۠Ox�LBd� �D$���q"����f$㛌�4�&F:pc��\�(�41b�x� u��A�b�����$�kB�Lj�,!	2c*|�h�?b2�%�͈��@�96)�c�/�bP�YoDnV�k��t���i" L� >�DS�a���%>�L~r���NBƳ���ĬeT�[b<��2�v6�Y(-��@BsN4�%�Q���H�b��М
�(5�Y@.>��N�c�%	O6��vA�N�&�y4�,�k�x�w�!L��( r�@'!�L�RЊ0SҠ���9��Ā�#	ѐ����8Gȁ�8Q��Xy�.Z��3!�IO��h>.(N�H���H��`s"����dr�1B�D������1�l<n��7��dd"2�)��2���1V���A ��qN�����s�(ޤLB:P'9�/Lh�d.E(A��4�q@]�n��9Qu�Ĥ�	�^�����H6��P���!0 2��d�C��Ü@̴�J`P���C�$ub�@"D�G&�X��Ar�Do� Ȉt&�J��31�1�p!8�d�cyb*������a(1�H\'��$nN�b<u��`� `H(I0��9
u��6M!b̀�@�7�|���h(���������Pȹ�V��b tC
�9 �PuC6 �H��5g1�3�~���ĸ�R���_
	'F��.>����t �:n��H@�u��g�Lf�rBAW0T�7Q�s�b�%��^�`~��i��N��C
�A"�N�eJbEp��T*��h(��/Jp�F»r;	�:u1`�20�t��d��tkE cC��1�|�1 "#0�Y|�QtC�uh!d���7TU�@H�f��R2r�e��
�
J|�>��c��e6��,XN��j0mo鶴i��v���ʃG����67qӢ f!NB�0�0&��N�е����ט�(��3��cق b� &5��A3��6uvѴ9�%c23s�v�L'�>g�Ԉ�956�UV�����_[UUU��D��s(�H]MW@ȍ �p���X�SW6VDCX�i'$�¨�Pv�g����,���H��Mb��,8�P(�~��?>���=��pH�r��&8L(�<a��K/7%�� �L�0�'#H\RҬ#n�s�9��xm'k�,���ov�2fL���/Ȫ<p��=�]~M	���[�@Ry�e��I��0,*�&-q H鹮��看�,O�vZ�4�}@D.�cRE�9g���iPU�����  Ǆa@*/]��>F���|���8B�f�����1�"��Sɖ��vޢY�}ǎ�X<!�[�t�D�&�,abw����lnGFs��㞳�
=D�jn��Py�q����B!H�΁�E���3�|�e�Ô��39F(\3��3	�-���,��,��  Il��q�#��|�%��Nfl� !C ���r�L�s-f�\r&�������,X8i�6rT���شqw<G4�d	Oy$@�*J��p"J�w	��pD"�F���������,X8e�S��W�㏶�Mb[�%�ߘ�g�c������y��y��3,9f�B�L���W̛?��Ӎ�1��&\��t	&B��%��*���-X�Eyt:m?����U ����䬋�qg�X�H�����D ˮh�B����#���BE�z�Ƞ��0��`粝]����2 QF��I�3͕جc���vCV��V�����s�yg?"D&��L.K���|��?�v��c�d�iRE�ed���9!.�@��}��SNi _�i���]�}'̺� ��,�
]�u]�4����	||?_Y.�CU��?���]�_fzZ%�u��1dZ��_ňA/�9�N]�UU������Y��a�`���A�g?j��k���q�]����)Q�\�3B"$n+����͡�;�,�2�@�tU�'UF��>y�sY�i(��01�����~�D�֏�����sΙ��ՃH�k`�yF���e��_�	9<�U�����ڀ:��eY>p�u} ��k��?9s��r8l��Nv��]�a!3�USg :�>}���eŀǽ�8�Zҏ�β,+��\p"US����`��I�iqؓs����1%�eFx8N.�R4"=I�`"����:O�է�,í.R�'N���ieP~avQQng�E ����PM�ҳ�i�d����2�upB�t�ea89�s��{��S� cX1elׄ�2 g��s��Q�4���V���k�MMM+W��eY��{�08�=�'���5�<X��GM�2y�̙�ON��ea� ��C��^�1ɲ�U^^�ĉSV�;G�*2c�! �h����{ҜgR4�=�cUU[[[���^xa��=��nw$ٵk�M7ߜ�����n�ۻ%R�4��W���������{���W�\�s������ҒҜ���f��̤Y0|��>X�r��,Y2޼���>ˊ��55��/,}aΜ9iiiD���'I� ��ZjIi> 0q�E�7C��Y�	�˲�ky*ܪU��~���Ɔ���{�g�9UUU������/#=��+�x�UW�l�S�!����=���h��g�}��7m�-Ѯ]���NM�f͜���}���v�d=�ea�����ƛo���+�f�l��}��t����|`B���"��o���+/��PUU״�/��}�������:k�--�F�Y Dٌ�l�$ BEa�ĒY�4�_X��ĉ����!�M�6���˅w�q��f[�v�+���x�⌌�n_����f�,˒�kzD����*Uw��`�AM��T2'Q��a�f}��+V̟?���
�~���|�fM/4�^��R��M��.]�d��sf�~����k�����?WL������D$"��iơF d"����A�K�����E�466�?~�ȑo�����W���v�����OgefN�1���E�n������UMmm]}= ̟7����ɏ��#_v�e�,7��TUUuk#�,�,��hw�ߟ���v�����Ng �\�{Y˖-U6����x<�)�.�� ?��_��V�X9����f�!03��HU�fn��T<C�����n��m�-^�x߾}?��+�vUֵ"�-������Ç炳�|>Q��.\�~������GyD\|Y��`�ͷ�
����ޮ�;��������?\�pᐍ  8p�����e�� w�uWJ� JJJ���<8���˽r"��Ed��yuΉ@�;St�����`�}O<�D<������;::~��C�s�К�1�4ztYWmHFb��b"�>�Y�.lUFFƬ�3����s����q�Ǝ5�o����gώF������ TU���[[[G����0%%e�ʲ0$㻧_i���O���r�  ��1c�o���NX���444�;f�e��|@H3Mi �d��tI�ڪ$��x��r�}��o��|��mӧM��k322*++%I궭{9��KYEEEy�y �v�����ѣG;v������gdd���tk��N���h6�At{�Hư������>��3�\�dIzz���G��߿��1i���(�;�v�dS���JI��=�ѣ�>��Ö��1 QZ
 /��2 ��,))�� �K5z*K�4MS%IR���V(N�K�T"RU��p��,)+�~zh�KYӦN����}�ٝ;w�1BU�={� �w|��v�ff�S  ���j&�b(�w&W=�X�[߼���.ݼi?���w|��*r��Z�,��q�7͜93/?��g�]�bEy����{oCCCiiiO��!?�k!I0�z��HO�8qb0<�zVVV�c e9��+�XR6�lժU��m,���srrz�IV�:��^��\hP��N��z�'�����x�	q1T�qEQzw��Vq���ʏ>Z=e��3f�,�"��`e�$I��3�����n�9�:$���̴Ȼd�4�w&�<cH:�$��T!6�z?]VVVVV6��,�	�'�d ���i+K��3f:9���E�|����,Ɉl(� �QeY>H�Ę44��k<aY�{؅j�3"Z!7q�s���,�,�r:˲0�L�ژ1�����?me�H�ľѮt�̀ ã�v_IJ^��β,�!eY��G�dYI�,v��꺜J0��Q@D&z��?��I���J�$�s�`�$���)��p2m���1�����Y��4#����O#�D��Q����V�$Ƙ��aʒ< �dIfȒ?�:�,7�E�u]�z2*"J�$Il ���,#裙F@F$�y2.6�j8d�(˜s]�-���� w���}��٠˲0|@DY��c�1Z��P��Q0B�^	�D�\BNH����PM�̸���Dd�0��OgY��"�$�I�ܤ�J�3��N���,4F d��5ߐw�4x�RN�R�t�ea��R:]�8�e����P$@��C�"�E2�h��5Λ1s�&$��cY�0���IF#1��K�\���`� �&�lxW���H�������D�
�F�3�����2�`a�f��H�GH��ryZ�`a���� 2�q�Sl9��;V#Y�0X��#�#q�L�:f	3�4�J!!d��H�K L��,X$��9M�;>!#�Hr �Xf� �(ƛ���h$�e$��,X�0� "���N�q������B�ׯ������6�C�'jnn~���+++UU+))���EEEE����xyF �� �t�����9VYY�ʫ�~��{�~����������#����;���?��������+����x�    IDAT�=��p�
�.g�e  Ƒ�{�p������G��'D\�n�O>y�ܳn��f��{��5k��������C��ҥ/�x��_�%�>�¬s��#.l��s�@�FΩ��n��m<�-�����M�w��w��C6�~�?�����A�r�0���ڲ}��Y���h �"HK\��1������կw�ڕ���/]���>�ֶ�t��hz9�w����(�� �q�l�������x�^K��������r�H2D���O3�􁋜�]]D�;w��z���ǟx��w��i�i���ݞ��� |���{��k�Q��w)��$9t	 4M������L</F$I"�Q�B@F�rb_� 8����{Y���3ft�.����G� ��9��K��$��EzR����4�0`i�W���e�j#��$ ���G<�i���\qŒի?nkkSU �N�Z1y����s����BWkh��}�Pu`���`�F��c������1c����A�/�Y/���i����0/���!��_p8��������K_| �|�M�7���{ǎ�;� �˲���}9&�|͌)k֮ ���3f��-��������p	!D�2��ӌ�k����3�.��B]�z��Ç[�ݛ0��n������_y�ޯ�rKff��J�_�4��R@�"F#��qYSf�,���n�5s&"Μ9s���6lضu[/�- @vv�̙3��P0ء�"�|�Y�f�{�S�N�f�;���������"��olh�;ש(��_ ��}�����V�����{﹧������s=��]V֋����3�B�	��H �HĹ�w�J*))�V�p*�N�I��v�?�$�2 b̈l��8��)�H�04�k>�q�SD���X�0"͈ ������<Gm���AA>D4NO���H�-X�0�ř����0 ��
�H@A,�,���Cx�d���o-�,X��\�2 ���B$ �-�т���3Ӛ�!!��Vh+K2C#D�	���X�Y�|�4v�	��Ȁ,{�C�2&�U��A#�;!�D�!�H��:qk˻�i	
�m�P�x��9������n�B�� K��eC��BSc�`��@�WD���vEL�-5��:m_�v����)�Y�Cw��80'�2��BeZ����U�=���Z��q��UoST%n�B��퐗ʊ}Ҵ"yJ����{4B8�#ʄ	�! 7�2�k��^��]��V�&�\�:���%{��U���4v���QJ�c���q8x\qslg���V/$�h䏀?��k��T�9^vI����T��!�!�dS��V�*Κ�|�����QU�zm�����q�w�W�Wn_��%����Z�;���hGԢ� Q��U�˚�Ǖ�W�:��8 ��Mi b	�"G B�4�����E^��86$��G�ߏ�<��Kَ���5��6Xp�]u�#D>9�@#@#�>"26��}�9��"���׭�2�i�����z-y9���wv�#��C��6��+«��M3�D �g\8�#A��Q�^��R�Y]2�h
��?�6�v������b�У=B�����5J��� I:7�����,6�j˶�-96L�vT{qK,��Ѽ����>�Zrl�d�??�c�i^d��8 "����Io��4zqs���a]��گֶ�6��:��%�Y�0\ �Ϫ՝u�Q�	��0� 1�C�4n:�U6�m��W�sa�SA X�7�؇���6��R�x����eC�[j�kz_�Hs���/�r�t��mkm�#��K|���[�Q�A��G��]�#�<+��O�����I:\�u����=��R��l��&�u�u�H��\%�I���@�����s�ψ�����G�
��h��;��/��o׶����0������Ӱ�TQh��´��|�/�'���n�M;v+�vӚC�rf���	�L����n�:��8]�D�a��6~�E��������ԫ}�_�P���2eCM'(��g����5|fN��Vk�(%�����KP8p@�rI�䴇��f=�ǻ2�z��iL�r�h��s��JY�쵳SKd��'�O�/��Rd�+��f��ֈ�2����q_���H�΅���侶��~��!����O��l�n�-�y�w���������r������<��§H ��rO*�;̵]�^��x�3�v�Th��}� �>�ֳ��u��i�+i���X� ���8pF �A���?B���&�]u�7����X{kG��{��~c[x��Ms=���kB�EUJq�@���xc@_�7�9��d�G�(���X��3wT^��x��#�wS#q>��&1�X���\l[m��Q�栞�*����#qU'����Ӝ,�+��y�0��V��[���ڸ�i�X��T�o��k�6����C+�߿�:?���z1�[�Ʌ�$���P��w/�r�wr��O�zud�<�ؖ�Z��[k���?��K�\6�G�Ks������`f�}�X[�W�����}����<ej�ݩ�?B��:�(�ex��mھ5�L.���m!}�1U�4��^Qh��µrOD�SKlN�nR�5�g��5�g�LJo��?�,����PO�s8�Q�۠23{�I�����3=�w�?�ML�:�c��i�Q�JL��� ��v�e��y׿�A����q�J �Gf��3�i%��T�8]~zC�-��]n������T5k߿(�!�3�4����[�Į��b��9�Gfɛ�c 0��q�|okH�K���$���hק~��mkM|HfG�L�mA����{�=	%�Sk�z�U�o���9w��Ǘ�yx�8G J����T�ˋ'8g��m��c�/�I��\�r���!|�l�/���ح�-!=/Uzb}�\6�K�K3�O�u3�Lt�c��������ѳ���Z����)�k[Con�J6��*���C���x�\�5����������p���Z42���ET(��z��C�WC�w��A����w�࿖�W�� LN_F�kO6?�>�tc��}��ܧ!���(��f�sG�^��+m����wv��z����/Mw��UDb������z�E�Qb��J�;_���ٖU{� �u�K+\�(_�#�����p�0�TM�>`��;�����[C��������s��=�bI(2��՟�ѦH�H��۾�@D�A&�I�q�Hcs�%=V6��.���G���� �;Ҿ�H�h��ޞ������]O�~����Gb���x캙�5#�x����/Lq�e�`_�5�?�~@Ȯ�F�}��go�ylt�r�I�H��$C ��� ��!CL�y�!0���桕��'9���\qBV�K�]%�W��}�U�0�I���S�3J�U�8�M���#�-��D�����9���k;��p�4�S$NQn��cG"�o�(� �	l2�I��cGZ4M�|*���[<H�vdy�O��#��)Q��k_B�	�Lv�:�d�d�k������c�dz�/��;��ӪX�u}׏W$��P�&}V�jִ.��ʡ5��5��|�mG���:Զj�IO�Pt��C\�d��4��ܟO2W_(�#H�	�d���
z�g��X���p�M;Ԥ����y���5NG۴���
���Y#�ڦ��eN �k�=6��~�Q��Ky�P����*g��<��Bq>>�>>O�K�N� ��Q�f�pk���$M�`�iէI���"q
�h�6�%_����|����}�x/w�����\x���/��Y��#�� p����	��/����7ۺ���v��*���&aKPF�4�	�661�U�ӆ�(i�&(�Ģq
�H�)�"��ᑚ:�i��4�ȶ�X<�M|^�cO�z�XGU��s1Fg+�.F �3�nL�c�	jF�(#����!Y�3z-���.�p��أ7d��5�T|)�ܱ�B������d����Hlv���R��!���=|�t׍s<b=��'�䲴�T��O��Fk�$?�4-���D��7���ؾwQ�]FMU�e[C��/J�΢����a����_[��p8�׏{� �d�Oe=�*/���i�b�~�}����)�Q�R]�փX�=��?W�ݻ8�9���= [j��s椰�"���\0��	T�^�j�\���E)ӊm�N��a�q�;���sF�pq��ы���8=�Y0�#�����,�A�n��֫w.��*���'�K2�g(�� ���"ѭ8 qιz�&}������������U�{4����T��~�y�� ��^��<#|�?��?њ䴡��ZB��:��t���P0��t�I�!�S�L�@Dq�1��8�MƸF��9H|.IbUI��=̳�R[��5Js1��?�e�n	�*1!���#���J�)'?5��Vl��ei�E���������G���x�������E^�Kҫ��o�z�@���
�����F�7s(���k����G���q`L%E���k��`.;r1��]�4�tjs�0��d	B1
Ƹ�
�s1��Q�Q.JOq0��?}.��b��uD��`$1x�oaZ�L;r�i��� %�@f9C������O�ۆ������<��#\�,��2���T	 B1��S���w^m�bn���p�1��J'n;u���/&Ԥ�-[�p���;��#��S�DS��̆��;�ڊ�+e{Y�.��/��;H��KS���A}t����{�IK����'L�12h���Dy z����4r�Nj|�n��D;s��3�HUY�T�������	�d�81"2S��#꼑����X{�-��e�; U��?�w��i��T�����_ۦ%Y}��M�-<ŤyD���hRo�ɲ�p�'�`�����	A" ��e�ځ�ȁI��_z�'����{w�n�e7�V��k�e�(�<��El���j�]�iIp�$�5IbR�����)b�1q��1 $[i�:ֹp�RQ [�0l�-vE��ӗ�������o��T��)����BB �P�� ����_ �L��l��l��!�ۆ��wL-�{�Ρ�78�[���á��g��)�wv�̈!q� �y©�?�-}}�#�c�J�lx�t����n'��;�v�Y�0�K�K�m_��ߏI#"������)��_��Y���e��Ųd��P��r���EΛf9l��OeY�/���)6K��^�p���9����u(�U"�;��	��h�9qab���Ů����߫Z��AL�x�h��I���t�Ȑ�=����؛���V���!�.����V$���ġ2_֍�	+>��B{�x�mg9./���+��Fk	�H�:qnE��GEp�Nȕ/�`�+9m?��s��3獵}x@��2�2�{[��k/�
�m86W�`�2�P�8s��dFH�Ŧ4"g$��6�ӥ;�vv��p�~����Ӭ��=�y�)N�Ma#2�l/k�,AA�q���)�#���Vn���<v�Ma%>V����fkz��i@"l�H�;$�ͼv�\(O.�z�_lG�+�ϵZ�tÌ� �DdoB�LDAE"��_,XE�䚌 ��/�D�iDn͂���3aR�	�ZMb�����dh�7CB��`��Dd�HV�i��k $�!Mk�[�):p+/�C�31
H&��u9��.�)�&'��޲L�;e��2���8�T�I ��9�� ��Yֿ�z-B��Q8Nq�t�3�WV��� >��Aj`�8�b�E��ƵA���s�I��!�(�;�D~��1�ƿ��N{���5�����V�=LQ�ڞ�"�tn
+N7rO�6��a�  �7�U  �u�C0]׉��U�> ����(ɒ�؀������[b;�V+�t��f��ߨ��T����i�ANz�277��xjbaF+��\׭ù�մ5U�I�<�����vŞ�Zy���JGZ������To��>���b�$B"U9F� 8���iǆ
�sM�8�����k"Ojql(���=�~ �����qE�ic�Ƒ#�����;&,�Ѫ�k��|��#���w���C��6����;e�)��02�DB$6 }]�-�� �B7������Xz�G��=md^Bd��e&B�˱o6�3�O{L�y5Y���5m�?��+�tgbid:u.��U9b�5�Xf�������X8nql��
��G��{��#������,�I[9�ԗ�HD�P����1I��^oJJJ"d��d�L�uY�1*��m[_��S�l~��1��%�����vG*�~e�@����$a���z��C���y���Z�|�iCz !�H@Fh� ��q~�'���۶-k��={Z[Z�رc�>{��E��I7���[��~Ƙ/�7mڴ���S_�k��#�G.����Ӹ��mܴ	�̙�U����drO����NY<���:�Ov�'����|���O2�-�$���"f�ˆg�q�#��C��|��bۇ��K&���W�|B�2!����P�̐��s�8����fz��h��&��3�<�F?���QJM"�v����)N�  ���$Ug"��{7�|��G�<��Ǐ_s��s�ι������O=��O�b���mٲ�>��ȑ#�?�����n9�cǎ��x㴵��i�֮[�n���t�)Q������0e���p�C�Ӈ���޺|G�ڙ�sǞ�k��r�SJ3�9:G��e Hs��يS���ʩ���l��tw�r���fy�.G���<o� ʲ�)'E��H��᫞|�i4���@@��:E$�dg��֪������w�y�MQ��g/8��/~q����|�ɂ��K/��$�q޼�����^z魷ފ�b�$m߾�����vO�0!###Aપ��UUD4f����Ҏ���۷{���Ǐ���VTT ���U�U"�ѣˊ����[��ݣi�������v����UU��ҒC�쬬)S�H��m��ZZ[232���fZ�������`c@|]G�G�z�{�xӉ�:�S�K'��7��
W�ۈ��iU,�����k:W`r�Mah�A�\��7�Ч��#qj	�w��p\f���p^��j�􆎎g#3���JsP�8���xKP�N���m�]u��3B��ߨ�K.�7��#�D]l H@«8�ua�\�v��n���k�O4��f�]p���[��Y�v���>���#���V�\�}ǎiӦ;�`0��3�8�cuu3�O���o$�����>z�X{{{jJ�]wݥi��?����u����_������].�/�'�Rzz�c�=��ѡ��{+V���X�f�G�?v�\�&��w�yW������kΜ��>�ܺu�|>_UU�9g�}&�»��}垞?�{-'�ћ;B��*��'�D�c�ڌ[N���DJ�+&����Dy�W�纎����w�=�����m�d�w����H,��ׁ.Geɧ,���an���Q}d�?�+ݻ8Uf  �.��l�8�sA�ێv/�9�}��Lp}N>�4!���,�.0�AgB�ġ��g�~6u�Ԃ�| X�v- lذ��sϱ�l�/Xt������'Ѭ��ZӴ`G���c���7n�~��c��6l�d���|�M�6EQ����>|����?��СC%%Ś����Ȳ��_�j��]m��c��^�`�رcw�ٳcǎk��&������� �KK��o�����G�y���^X�~��#G|���n�����{��G��{�_﹧{�t�I�إSc}n���8�˳=��G�>�t7��T�+�C˶��y������;� �ܡ�狭��f�ۮ�7��F5��ڠ�ӁFgK����S��������v�,wn�|�(��ͮ�kSy��Ë� `r������'A�����K�������{�:��!!"gd�G���t(v�\�� ���} ��l�4������5���#�h��?��O����c�6mloo��׭_��iZg�h4��sϽ�lY8"MS %�y�^����srr�������z��7�x#��Q[[��n����RRR ��r���p�X1�  �IDAT׬Y�؟�r��I��X<�(6%++m�팠YϊC����=[R�qROQ�b*k{x�D�co�I�KB������u����(`�P$�����ޫ{���� �r��@b K��b���NU�>v(� Q��O��3���?�Q)��0$`DɐbDDdX��������܆��H8 �\}�����m�q������ݛ�K��OMt���oj"���Ԫ��ښ�ɓ'�/b����Ç��l�2j���I����������rˤI�v�ޝ�����Ș7o�̙3SSS�޹u�6��3fx� ���B��[�:|����g�0롩��R|r8ړI��rWM�V�ލ��R�X[�'�H���c*�e���a�]?U���?�猴/�D�H���R~Z�<�s�8ظ<e\���X�@�
 �ñ6}L�R�o��[U�F �}���'����A�LOR2�ˉ#D ��HX������d�O�cR�r��9�=��᪪I��eee?��O ::v��5~������Y�j�֭[u]///�?>�|�g�~&==]`��QD�v�ڱcǾ�λ���I��w[z[[�c������W^Y6jԵ�^��U>ݐ�����0q��(O=��c��h,�������dɒ�^{m���Lb�$�4뾃E��^��*c�-Zi�	$�0{��I�ww���.�4zp�_�����s=��A������N��`t��Ms܇��kF�yn��g{��_��-5�����#mӯ��o7�ꬭ�N)�����@M����K+\�u���O_o;NV��'5�Ѹ�J��/�[@2���9�.�x�O/��H�����z���~�;I�~s��]�f�>���+����Ӧu=---���$In���t����bv�]�4���9����,˲
�E �á(Jkkkzz:c�����p��v�߯i�,�^�WQUU;�A]�EIMM�����|�"�@@������+�b �d�N��t��(���g�iD�3�q��)#�8Ԥ>�n��2�	�=u�_����Ѓ>7�u�J���#\b��d���8�b��8�̌<�n�쬩C�:�ӆ�a�9�� ���-��>7�	�
�5b�q�ؙˆ�
l��������6	��%�k�vde�<}��ϼ���i�����Sd C3J�P%#��Ě�w0�z�Yvv�7o����("&�U�8m�Բ���8 	{}Wt��D����n�Iŉ���O�!!�һX\�^o�_�T��W��`=�V$�T�[�i"�p8�ү��(����ɨj�^�\�#|� ��ĝnHd���ə���r�8��:�������q�33u �y=�Ŧ��U��s4��:�&nn	�A��eYR~r��[Z� d(�(�@�` 90����NwR4�J�S1jԨQ�F�tq	`�?6F֫�Z�/�̔���{��5��{ϟ�fN9A �[C�v����8��V��4���>
��N!���NL*H"VW5�"ȝ��D�� ��
���d�(I���,�(c�W?�T'~i�}W_��C1�����o��ɽ0)_����4���5�N@�ŊB�q��$�Q3�,?�a�|H��g_�,��e�.8�jj���UU߿�:73C��0L�q����U'ID�d��ô얥d:¡�7�;��X����c_�e�?*��ӈ�{Wucc"
	Đ1����$1 ���u��gC�e,�9�$Ib��%��;X������޾�2�6ӗ!���;=�����M{���S���PWT��3f�bT���+�g[���� ��n�］?����BkV�ǴN}iT�����0@�$�p�tۧ����R���w����W�yֻ�d���9�MoN.�Z%Q�E���O~�'?�O(��P�R�@m����F;[	��	��If1f��"���4���z���z�}Nb�E���~ə�o��^�<�Y�����f�zM�6m]�Ϻ�����n;��.������^F��Ӈ�w���d�]�R�y�����_�~k/��  ��-?��CL��I,/_�z���8~�[�Ic̬�~�	۷of�l��6MSk��\���~���;[�o�+��V��ڟ���j�ᦣܾ�~�������9z筭]����o~��G��Lt�aF4M,�/g	Fn����_����=?����4M�kg�oCb����p2���~�����#ϼ<���u��/��=}�zgO�|�����W��`H�鲩7ԯ��D�,�Ճ����?t���u��wPi�뺯u����u������x�j��9F�$̄���y���F�C�v�����\�[��^��F����}��}YRN��`�I�db�'#)
x쑧N~����z�� ������J�P�q�DW6nT�%h�q�����o?|��&W�~���ul�.���ܹ�FS���O�Q爵.T�d�E��{y����_��ji�^��lo��7>�G��S���F���l���(�QQ4F��ړE�x���=w�����Λ���z�Wı�~��ɧOn63وA���(��۾�^$z�$���U�9z��+O<~�VK[��"y���_��O���~!l,HE��. mg��b�p��$#oEd�(���<efw��m��
 ��Mz����g�#p�o��߀FXD���,Z1���{�o,�D��f��V���+�>��/���ַ�|�֛֝���
bf�W�>��ÿ���Ϗ?�B�X�0�Pf6
�����s+8�Q�D&	4�u*s:��'�?����ں�Ǐ]O��כ��؛��ُ�ʧ����x�B�Uj�Ժ�Ŭ@(������`DP�q	w����8J��\r�����������޻Nܹ=m�:�}����`$_z�©Sg���}�Ͼ����m�$E����A��ވ���o�~F}�$ R1�7�<�p9��=;cN��-���w~�m������[o䁡��խ��=�`���������'�ʗN�=��K�E�+c��_��8�L;����ḡ����H��Iy�3L�!8$̂ 9<vI����[�u�������M7~�7�bv��}�Z4wd~������GF�;�ثX�������FΉ<%~H�.�o���G�f`�����9�)��T�X/R�S<)�����#c�\�k:D.��|p�<(�CnO��0wA6	�΋�c#]9��r��=���{J��g��u��������e�(xA���}H(�?���_�����/=��KgϞ;��7.^���fEw�X+��@鋒ؗ/#ڔ53X.�!io����% 6P&A�c�+�9�⿝}�zs��A�+���(5����@�CH�3�|��F	��#���_�u�E�(�zܐ2Ŏu�^���)��9�cG��M�wgw}�0Dg��Q�.���U_�n;�JBe��,1�-����#�b��S��dTuk�0��QxNK(!e&�RHDlx�گ�3$����VyF����M��) 3��{3�9Ei��Y���tV|%�rh����5A}��(́�rB�I�����ds~mm�/bY�rg��Ӥ�Ut�Ŷ*
�2"��iV�u^�S=��� L L�O�BC�!�}X�\%#!������hh��V�@�A�R|ShK���- �\�|�C�Z�[ �0��X߰*ϼUP�&�K4�ŗ��s<a.�Ŧ%R�&F4�b����=���x0�J�Pbp`�Z��4b*N��@�7M�+1����Y��R�(��`/�bI&����r��$��"�H
�zI���p�(�7 -���J4dj{,$�;q'�=�p�.�%�#<��NN���T�@A|+-f����DY��&�� �}��N���3�7@���n��<Ѳ�	8Zx����/B�ӧP2PS��a�G~)�R�`|aU(��D7��1�Q�9a�I�e��J� y d�W021�vy�|�������7]d'�N8�f"�a�t[�I�&�X>�=!N�fn��`^�8V�v/�(��g�&��-1�e�4B��5X����0f�+�9#7��rE�v�	�ZTg+����.�k3"-���[�(A�%�DK��s N24���6I��B �݂��0G|-�$|��0o�gŇ�#h�@�4�
z/h��R�)�9��b=��@T&cK_�&�A�B����06���F�q�+S�t0C�0�,rG�a�0'(�h3�놑U������#�qf�<3��|f�	�W�F0$3�r�p*nz̔��汏-4��|��:�4�\ �d��D�B	���it�h�t����4��b��:��0��(� �eE��S)�����vi�;̀F6S�
EX��y�/��� -[d�4��T5�4������G��c�*O�0�4��t�'D�����'�iyV�*P]�cAe�b�{��D!ҩ�r8e��3<:3�R�� �b�dDƪ����HF�T�9�z�8t3�E�(��$4+��n�#D7	2��-�Q�@o����F���h��9Ѱ�����%EF����X��%���ob@������i��,[��p�s�0C�bT`��d����@U�5�� ��B.Ll�`�4Z�E�%扑��}�37���Oa�l�T\	G�l2����C$�2%,�5B��.ͳ��Ƣ��ᬍ(�$)�I�G{����YT��25.F����	�����
�`�A�IR'��N�8d#uAe9����9#�HA����C�og����e0�p��V'%Y�fW�Br���?3	+ᨣ��{f�V�K�
/*Q��Yx��D[�
��R)�0SOk�ޗ�!�<+�7J	���&KR	A����}�"Xͥ[�$a�^#(��)U��5Ʌ�L��3,�׌h"@4���E�$�r�	}O���B�J��0�g�gwyڵ֑ֆ@$u�e�)ޤ�´=�=b���TZŞNAk/Ѝ/�5���P2	KE�&P�9�$��)�ŧ;n�(UJ��h-+�"
q;c�" �c��X}�=ֹQ��3G��^"s�!���(�[���ɕ����H"���1��gT�������r�B�X=ܭ�����茟.�4�Irv�	^Tf_y%@��\4ި�>5$@�x<�i�N�z
7��@>�;�b�%b�n'V*7ʌ�)=�͛Y���R$J6|k�|��C�N���y����p��[�,�(�}/J+HRbk�����ɝ����A�җP��n1�s�}�tZ�C�oXU�c�ܑ���x��@�d��'KD��Q�_�>��(Ŕ�}����SF����d�	,��x��qY8�e6]�G��<؜��(O
���ٝ� 	�H]0�����T�:XVOzA�ީ�X?�:��6��t�q�GOع(�u�<L����H0�|Rⶀ�X-��� ���R�g�F󾰉=C]�0��DyF����쾿�yS���!;�Mt�L}��v���e�Bi���ͺKF]>`���J�Ƨ+�Q.((b��+5Z,/#%�u
�erG=��t`��q�9Yj�,����;k�eN�=<9ʤ�Q��eY��5�[I���k�8�� G�uE;Je�R���`� �r���ዔ׽�f�2à�e�L/	�`Tڠ�F<�j\8��j]e�@D��(''�����F��Ε [��r���� u��JfY,bp���#=СD���.��M���Yi�L��c��Y�獪V�e �"�F�4e�TU���8���p��0:��y�mu�$�ک ��H��{���h�)�qFA��m�hZ�l����;Gٻ��nf�M���2�E�ԣʣCӒ�����Q��z�2Du*��3,�w��yZ�ڹF�a�w�\��G�*� l��:��Lw�.����SU�YD���G��WTe�E���mhUz���Ի��3,��:Jԡ:��zb)P%R�E�E�,4�\��屺��jUG� A>C��hF���[/�͒���z݊*E	���o$Źd\T��Z�D�,�w0 �Wam�I)��ap}OE�DZ���G�40�@.����𖥸�    IEND�B`�