<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Window operations</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Desktop</a> › <a class="trail" href="shell-overview.html#apps" title="Program och fönster">Program och fönster</a> » <a class="trail" href="shell-windows.html" title="Fönster och arbetsytor">Fönster och arbetsytor</a> › <a class="trail" href="shell-windows.html#working-with-windows" title="Arbeta med fönster">Windows</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Window operations</span></h1></div>
<div class="region">
<div class="contents"><p class="p">Windows can be resized or concealed to suit workflow.</p></div>
<div id="min-rest-close" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Minimize, restore and close</span></h2></div>
<div class="region"><div class="contents">
<p class="p"> To minimize or hide a window:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Click the <span class="gui">-</span> in the top left hand corner of the application's <span class="gui">menu bar</span>. If the 
       application is maximized (taking up your whole screen), the menu bar will appear at the very top
       of the screen. Otherwise, the minimize button will appear at the top of the application window.</p></li>
<li class="list"><p class="p">Or press <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Space</kbd></span></span> to bring up the
       window menu.  Then press <span class="key"><kbd>n</kbd></span>. The window 'disappears' into the
       Launcher.</p></li>
</ul></div></div></div>
<p class="p">To restore the window:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list"><li class="list"><p class="p">Click on it in the <span class="link"><a href="unity-launcher-intro.html" title="Använda programstartaren">Launcher</a></span>
       or retrieve it from the window
       switcher by pressing <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Tab</kbd></span></span>.</p></li></ul></div></div></div>
<p class="p"> To close the window:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Click the <span class="gui">x</span> in the top left hand corner of the window, or</p></li>
<li class="list"><p class="p">Press <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F4</kbd></span></span>, or</p></li>
<li class="list"><p class="p">Press <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>Space</kbd></span></span> to bring up the
       window menu.  Then press <span class="key"><kbd>c</kbd></span>.</p></li>
</ul></div></div></div>
</div></div>
</div></div>
<div id="resize" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Resize</span></h2></div>
<div class="region"><div class="contents">
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">A window cannot be resized if it is <span class="em">maximized</span>.</p></div></div></div></div>
<p class="p">To resize your window horizontally and/or vertically:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list"><li class="list"><p class="p">Move the mouse pointer into any corner of the window until it changes into a
 'corner-pointer'. Click+hold+drag to resize the window in any direction.</p></li></ul></div></div></div>
<p class="p">To resize only in the horizontal direction:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list"><li class="list"><p class="p">Move the mouse pointer to either side of the window until it changes into a
 'side-pointer'.   Click+hold+drag to resize the window horizontally.</p></li></ul></div></div></div>
<p class="p">To resize only in the vertical direction:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list"><li class="list"><p class="p">Move the mouse pointer to the top or bottom of the window until it changes
 into a 'top-pointer' or 'bottom-pointer' respectively.   Click+hold+drag to
 resize the window vertically.</p></li></ul></div></div></div>
</div></div>
</div></div>
<div id="arrange" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Arranging windows in your workspace</span></h2></div>
<div class="region"><div class="contents">
<p class="p">To place two windows side by side:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Click on the <span class="gui">title bar</span> of a window and drag it toward the
  left edge of the screen.  When the <span class="gui">mouse pointer</span> touches the edge,
  the left half of the screen becomes highlighted. Release the mouse button and
  the window will fill the left half of the screen.</p></li>
<li class="list"><p class="p">Drag another window to the right side: when the right half of the
  screen is highlighted, release. Each of the two windows fills half the
  screen.</p></li>
</ul></div></div></div>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Pressing <span class="key"><kbd>Alt</kbd></span> + click anywhere in a window will allow you to
       move the window. Some people may find this easier than clicking on the
       <span class="gui">title bar</span> of an application.</p></div></div></div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-windows.html#working-with-windows" title="Arbeta med fönster">Arbeta med fönster</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links "><a href="unity-menubar-intro.html#window-management" title="Window management buttons">Window management buttons</a></li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
