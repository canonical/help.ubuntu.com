<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>What is the HUD?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Desktop</a> › <a class="trail" href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">What is the HUD?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">The <span class="gui">HUD</span> or <span class="gui">Heads Up Display</span> is a search-based 
alternative to traditional menus and was introduced in Ubuntu 12.04 
LTS.</p>
<p class="p">Some apps like <span class="link"><a href="https://apps.ubuntu.com/cat/applications/gimp" title="https://apps.ubuntu.com/cat/applications/gimp">Gimp</a></span> or 
<span class="link"><a href="https://apps.ubuntu.com/cat/applications/inkscape" title="https://apps.ubuntu.com/cat/applications/inkscape">Inkscape</a></span> have hundreds of menu items. If 
you're using apps like these, you may remember the name of a menu option, 
but you might not remember how to find it in the menus.</p>
<p class="p">Using a search box can be quite a bit faster than navigating extended 
menu hierarchies. The HUD also can be more accessible than normal menus as 
some people are unable to precisely control a mouse pointer.</p>
</div>
<div id="use-the-hud" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Use the HUD</span></h2></div>
<div class="region"><div class="contents">
<p class="p">To try the HUD:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Tap <span class="key"><kbd>Alt</kbd></span> to open the HUD.</p></li>
<li class="steps"><p class="p">Start typing.</p></li>
<li class="steps"><p class="p">When you see a result that you want to run, use the up and down 
      keys to select the result, then press <span class="key"><kbd>Enter</kbd></span>, or click 
      your desired search result.</p></li>
<li class="steps"><p class="p">If you change your mind and want to exit the HUD, tap the 
      <span class="key"><kbd>Alt</kbd></span> again or the <span class="key"><kbd>Esc</kbd></span>. You can also click 
      anywhere outside the HUD to close the HUD.</p></li>
</ol></div></div></div>
<p class="p">The HUD keeps track of your search history and adjusts the search 
results to be even more useful the more you use it.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
