<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Diskar och lagring</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Diskar och lagring</span></h1></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="linkdiv "><a class="linkdiv" href="disk-partitions.html" title="Hantera volymer och partitioner"><span class="title">Hantera volymer och partitioner</span><span class="linkdiv-dash"> — </span><span class="desc">Förstå vad volymer och partitioner är och använda diskverktyget för att hantera dem.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="disk-resize.html" title="Justera storleken på ett filsystem"><span class="title">Justera storleken på ett filsystem</span><span class="linkdiv-dash"> — </span><span class="desc">Förminska eller förstora ett filsystem och dess partition.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="disk-check.html" title="Kontrollera din hårddisk efter problem"><span class="title">Kontrollera din hårddisk efter problem</span><span class="linkdiv-dash"> — </span><span class="desc">Testa din hårddisk för att kontrollera att den är frisk och utan problem.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="disk-capacity.html" title="Kontrollera hur mycket diskutrymme som finns kvar"><span class="title">Kontrollera hur mycket diskutrymme som finns kvar</span><span class="linkdiv-dash"> — </span><span class="desc">Använd <span class="gui">Diskanvändningsanalysatorn</span> eller <span class="gui">Systemövervakaren</span> för att kontrollera utrymme och kapacitet.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="disk-repair.html" title="Reparera ett skadat filsystem"><span class="title">Reparera ett skadat filsystem</span><span class="linkdiv-dash"> — </span><span class="desc">Kontrollera om ett filsystem är skadat och för tillbaka det till ett användbart tillstånd.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="addremove-creator.html" title="Skapa en startdisk"><span class="title">Skapa en startdisk</span><span class="linkdiv-dash"> — </span><span class="desc">Konvertera ett USB-minne till en enhet från vilken du kan starta och installera Ubuntu.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="disk-format.html" title="Ta bort allt från en flyttbar disk"><span class="title">Ta bort allt från en flyttbar disk</span><span class="linkdiv-dash"> — </span><span class="desc">Ta bort alla filer och mappar från en extern hårddisk eller USB-enhet genom att formatera den.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="disk-benchmark.html" title="Testa din hårddisks prestanda"><span class="title">Testa din hårddisks prestanda</span><span class="linkdiv-dash"> — </span><span class="desc">Kör prestandatester på din hårddisk för att kontrollera hur snabb den är.</span></a></div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="hardware.html" title="Maskinvara och drivrutiner">Maskinvara och drivrutiner</a><span class="desc"> — <span class="link"><a href="hardware.html#problems" title="Vanliga problem">Hårdvaruproblem</a></span>, <span class="link"><a href="printing.html" title="Utskrifter">skrivare</a></span>, <span class="link"><a href="power.html" title="Ström och batteri">ströminställningar</a></span>, <span class="link"><a href="color.html" title="Färghantering">färghantering</a></span>, <span class="link"><a href="bluetooth.html" title="Bluetooth">Bluetooth</a></span>, <span class="link"><a href="disk.html" title="Diskar och lagring">diskar</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
