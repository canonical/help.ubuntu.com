<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Lägg till ett konto</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Inställningar</a> » <a class="trail" href="accounts.html" title="Nätkonton">Nätkonton</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Lägg till ett konto</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Att lägga till ett konto kommer att hjälpa dig att länka dina nätkonton med ditt GNOME-skrivbord. På så sätt kommer ditt e-postprogram, chattprogram och andra liknande program att ställas in åt dig.</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Nätkonton</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Nätkonton</span> för att öppna panelen.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">+</span>-knappen i nedre vänstra hörnet av fönstret.</p></li>
<li class="steps"><p class="p">Välj typen av konto som du vill lägga till.</p></li>
<li class="steps"><p class="p">Ett litet webbplatsfönster eller dialogruta kommer att öppnas där du kan mata in dina autentiseringsuppgifter för ditt nätkonto. Om du till exempel ska ställa in ett Google-konto så mata in ditt användarnamn och lösenord från Google. Vissa leverantörer låter dig skapa ett nytt konto från dialogrutan för inloggning.</p></li>
<li class="steps"><p class="p">Om du har matat in autentiseringsuppgifter korrekt så kommer du att bli tillfrågad om du vill ge GNOME behörighet att nå ditt nätkonto. Ge behörighet för att fortsätta.</p></li>
<li class="steps"><p class="p">Alla tjänster som erbjuds av en kontoleverantör kommer att vara aktiverade som standard. <span class="link"><a href="accounts-disable-service.html" title="Styr vilka nättjänster ett konto kan användas med">Slå om</a></span> individuella tjänster till <span class="gui">AV</span> för att inaktivera dem.</p></li>
</ol></div></div></div>
<p class="p">Efter att du har lagt till konton, kan program använda de kontona för de tjänster du har valt att tillåta. Se vidare i <span class="link"><a href="accounts-disable-service.html" title="Styr vilka nättjänster ett konto kan användas med">Styr vilka nättjänster ett konto kan användas med</a></span> för information om hur du styr vilka tjänster som ska tillåtas.</p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">Många nättjänster tillhandahåller ett autentiseringselement som GNOME sparar istället för ditt lösenord. Om du tar bort ett konto, bör du också återkalla det certifikatet i nättjänsten. Se <span class="link"><a href="accounts-remove.html" title="Ta bort ett konto">Ta bort ett konto</a></span> för vidare information.</p></div></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="accounts.html" title="Nätkonton">Nätkonton</a><span class="desc"> — <span class="link"><a href="accounts-add.html" title="Lägg till ett konto">Lägg till ett nätkonto</a></span>, <span class="link"><a href="accounts-remove.html" title="Ta bort ett konto">Ta bort ett konto</a></span>, <span class="link"><a href="accounts-which-application.html" title="Nättjänster och program">Lär dig om tjänster</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
