<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>The internet seems slow</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html" title="Nätverk, webb, e-post &amp; chatt">Nätverk, webb, e-post &amp; chatt</a> » <a class="trail" href="net-problem.html" title="Nätverksproblem">Nätverksproblem</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">The internet seems slow</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">If you are using the internet and it seems slow, there are a number of things that could be causing the slow down.</p>
<p class="p">Try closing your web browser and then re-opening it, and disconnecting from the internet and then reconnecting again. (Doing this resets a lot of things that might be causing the internet to run slowly.)</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list">
<p class="p"><span class="em-bold em">Busy time of day</span></p>
<p class="p">Internet service providers commonly setup internet connections so that they are shared between several households. Even though you connect separately, through your own phone line or cable connection, the connection to the rest of the internet at the telephone exchange might actually be shared. If this is the case and lots of your neighbors are using the internet at the same time as you, you might notice a slow-down. You're most likely to experience this at times when your neighbors are probably on the internet (in the evenings, for example).</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Downloading lots of things at once</span></p>
<p class="p">If you or someone else using your internet connection are downloading several files at once, or watching videos, the internet connection might not be fast enough to keep up with the demand. In this case, it will feel slower.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Unreliable connection</span></p>
<p class="p">Some internet connections are just unreliable, especially temporary ones or those in high demand areas. If you are in a busy coffee shop or a conference center, the internet connection might be too busy or simply unreliable.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Low wireless connection signal</span></p>
<p class="p">If you're connected to the internet by wireless (wifi), check the network menu on the menu bar to see if you have good wireless signal. If not, the internet may be slow because you don't have a very strong signal.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Using a slower mobile internet connection</span></p>
<p class="p">If you have a mobile internet connection and notice that it is slow, you may have moved into an area where signal reception is poor. When this happens, the internet connection will automatically switch from a fast "mobile broadband" connection like 3G to a more reliable, but slower, connection like GPRS.</p>
</li>
<li class="list">
<p class="p"><span class="em-bold em">Web browser has a problem</span></p>
<p class="p">Sometimes web browsers encounter a problem that makes them run slow. This could be for any number of reasons - you could have visited a website that the browser struggled to load, or you might have had the browser open for a long time, for example. Try closing all of the browser's windows and then opening the browser again to see if this makes a difference.</p>
</li>
</ul></div></div></div>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-problem.html" title="Nätverksproblem">Nätverksproblem</a><span class="desc"> — 
      <span class="link"><a href="net-wireless-troubleshooting.html" title="Wireless network troubleshooter">Troubleshooting wireless connections</a></span>,
      <span class="link"><a href="net-wireless-find.html" title="I can't see my wireless network in the list">finding your wifi network</a></span>…
        </span>
</li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
