<!DOCTYPE html>
<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Vad är överlagda rullningslister?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 16.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="shell-overview.html" title="Skrivbord, program &amp; fönster">Skrivbord</a> › <a class="trail" href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Vad är överlagda rullningslister?</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Ubuntu inkluderar <span class="em">överlagda rullningslister</span>, vilket tar upp mindre plats på skärmen än vanliga rullningslister och ger dig mer utrymme för det du jobbar med. Även om inspirationen kom från mobila enheter, där vanliga rullningslister inte behövs, är Ubuntus överlagda rullningslister utformade för att fungera lika bra med en mus.</p>
<p class="p">Vissa program som Firefox och LibreOffice har ännu inte stöd för de nya rullningslisterna.</p>
</div>
<div id="using" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Att använda rullningslisterna</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Den överlagda rullningslisten visas som en tunn orange remsa vid kanten av ytan som kan rullas. Rullningslistens position motsvarar skärmens position i det rullningsbara innehållet. Remsans längd motsvarar innehållets längd; ju kortare remsa, ju mer innehåll.</p>
<p class="p">Placera din muspekare över valfri punkt på den rullningsbara kanten av innehållet för att visa <span class="gui">tumreglaget</span>.</p>
<div class="list"><div class="inner">
<div class="title title-list"><h3><span class="title">Sätt att använda rullningslisterna:</span></h3></div>
<div class="region"><ul class="list">
<li class="list"><p class="p">Dra <span class="gui">tumreglaget</span> upp eller ner för att flytta skärmens position exakt dit där du vill ha den.</p></li>
<li class="list"><p class="p">Klicka på rullningslisten för att flytta skärmens position exakt dit där du vill ha den.</p></li>
</ul></div>
</div></div>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="shell-overview.html#desktop" title="Skrivbordet">Skrivbordet</a></li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="mouse-touchpad-click.html" title="Klicka, dra eller rulla med styrplattan">Klicka, dra eller rulla med styrplattan</a><span class="desc"> — Klicka, dra eller rulla via tryckningar och gester på din styrplatta.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
