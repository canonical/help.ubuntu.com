<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Mata in speciella tecken</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="tips.html" title="Tips och tricks">Tips och tricks</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Mata in speciella tecken</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan mata in och titta på tusentals tecken från de flesta av världens skriftsystem, till och med de som inte finns på ditt tangentbord. Denna sida listar några olika sätt på vilka du kan mata in specialtecken.</p>
<div role="navigation" class="links sectionlinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Metoder att mata in tecken</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="tips-specialchars.html#characters" title="Tecken">Tecken</a></li>
<li class="links "><a href="tips-specialchars.html#compose" title="Compose-tangent">Compose-tangent</a></li>
<li class="links "><a href="tips-specialchars.html#ctrlshiftu" title="Kodpunkter">Kodpunkter</a></li>
<li class="links "><a href="tips-specialchars.html#layout" title="Tangentbordslayouter">Tangentbordslayouter</a></li>
<li class="links "><a href="tips-specialchars.html#im" title="Inmatningsmetoder">Inmatningsmetoder</a></li>
</ul></div>
</div></div>
</div>
<div id="characters" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Tecken</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Ett annat användbart program som följer med GNOME är <span class="app">Tecken</span>. Det låter dig söka efter och infoga ovanliga tecken genom att bläddra genom teckenkategorier eller leta efter nyckelord.</p>
<p class="p">Du kan starta <span class="app">Tecken</span> i översiktsvyn <span class="gui">Aktiviteter</span>. För mer information om Tecken, se <span class="link"><a href="help:gnome-characters" title="help:gnome-characters">handboken för Tecken</a></span>.</p>
</div></div>
</div></div>
<div id="compose" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Compose-tangent</span></h2></div>
<div class="region"><div class="contents">
<p class="p">En Compose-tangent är en speciell tangent som låter dig trycka ner flera tangenter i rad för att få ett specialtecken. För att till exempel skriva det apostroferade tecknet <span class="em">é</span> kan du trycka på <span class="key"><kbd>compose</kbd></span> och sedan <span class="key"><kbd>'</kbd></span> och sedan <span class="key"><kbd>e</kbd></span>.</p>
<p class="p">Tangentbord har inte specifika compose-tangenter. Istället kan du definiera en av de existerande tangenterna på ditt tangentbord som en compose-tangent.</p>
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">Du måste ha <span class="app">Justering</span> installerat på din dator för att ändra denna inställning.</p></div></div></div></div>
<div class="steps"><div class="inner">
<div class="title title-steps"><h3><span class="title">Definiera en compose-tangent</span></h3></div>
<div class="region"><ol class="steps">
<li class="steps"><p class="p">Öppna översiktsvyn <span class="gui"><a href="shell-introduction.html#activities" title="Översiktsvyn Aktiviteter">Aktiviteter</a></span> och börja skriv <span class="gui">Justering</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Justering</span> för att öppna programmet.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Tangentbord &amp; mus</span>-fliken.</p></li>
<li class="steps"><p class="p">Tryck på <span class="gui">Inaktiverad</span> intill inställningen <span class="gui">Compose-tangent</span>.</p></li>
<li class="steps"><p class="p">Slå på växeln i dialogen och välj tangentbordsgenvägen du vill använda.</p></li>
<li class="steps"><p class="p">Kryssa i kryssrutan för den knapp du vill använda som Compose-tangent.</p></li>
<li class="steps"><p class="p">Stäng dialogrutan.</p></li>
<li class="steps"><p class="p">Stäng fönstret <span class="gui">Justering</span>.</p></li>
</ol></div>
</div></div>
<p class="p">Du kan mata in många vanliga tecken genom att använda compose-tangenten, till exempel:</p>
<div class="list"><div class="inner"><div class="region"><ul class="list">
<li class="list"><p class="p">Tryck <span class="key"><kbd>compose</kbd></span> sedan <span class="key"><kbd>'</kbd></span> och sedan ett tecken för att placera en akut accent ovanför det tecknet, som till exempel <span class="em">é</span>.</p></li>
<li class="list"><p class="p">Tryck <span class="key"><kbd>compose</kbd></span> sedan <span class="key"><kbd>`</kbd></span> och sedan ett tecken för att placera en grav accent ovanför det tecknet, som till exempel <span class="em">è</span>.</p></li>
<li class="list"><p class="p">Tryck <span class="key"><kbd>compose</kbd></span> sedan <span class="key"><kbd>"</kbd></span> och sedan ett tecken för att placera ett trema ovanför det tecknet, som till exempel <span class="em">ë</span>.</p></li>
<li class="list"><p class="p">Tryck <span class="key"><kbd>compose</kbd></span> sedan <span class="key"><kbd>-</kbd></span> och sedan ett tecken för att placera ett makron ovanför det tecknet, som till exempel <span class="em">ē</span>.</p></li>
</ul></div></div></div>
<p class="p">För ytterligare compose-tangentsekvenser se <span class="link"><a href="http://en.wikipedia.org/wiki/Compose_key#Common_compose_combinations" title="http://en.wikipedia.org/wiki/Compose_key#Common_compose_combinations">compose-tangentsidan på Wikipedia</a></span>.</p>
</div></div>
</div></div>
<div id="ctrlshiftu" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Kodpunkter</span></h2></div>
<div class="region"><div class="contents">
<p class="p">Du kan mata in vilket Unicode-tecken som helst genom att använd bara ditt tangentbord med tecknets numeriska kodpunkt. Varje tecken identifieras med en fyra-teckens kodpunkt. För att hitta kodpunkten för ett tecken, hitta tecknet i teckentabellprogrammet och titta i statusraden eller fliken <span class="gui">Teckendetaljer</span>. Kodpunkten är de fyra tecknen efter <span class="gui">U+</span>.</p>
<p class="p">För att mata in ett tecken via dess kodpunkt, håll ner <span class="key"><kbd>Ctrl</kbd></span> och <span class="key"><kbd>Skift</kbd></span> och skriv <span class="key"><kbd>U</kbd></span> följt av den fyra tecken långa kodpunkten, och släpp sedan <span class="key"><kbd>Ctrl</kbd></span> och <span class="key"><kbd>Skift</kbd></span>. Om du ofta använder tecken som du inte kan nå enkelt med andra metoder kan det vara värdefullt att memorera kodpunkterna för de tecknen så att du kan mata in dem snabbt.</p>
</div></div>
</div></div>
<div id="layout" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Tangentbordslayouter</span></h2></div>
<div class="region"><div class="contents"><p class="p">Du kan få ditt tangentbord att bete sig som ett tangentbord för ett annat språk, oavsett vilka tecken som finns tryckta på tangenterna. Du kan till och med enkelt byta mellan olika tangentbordslayouter via en ikon på systemraden. För att lära dig hur, se <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa tangentbordslayouter">Använd alternativa tangentbordslayouter</a></span>.</p></div></div>
</div></div>
<div id="im" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Inmatningsmetoder</span></h2></div>
<div class="region"><div class="contents">
<p class="p">En inmatningsmetod expanderar de föregående metoderna genom att tillåta inmatning av tecken inte enbart med tangentbordet utan också andra inmatningsenheter. Du kan till exempel mata in tecken med en mus via en gestmetod eller mata in japanska tecken via ett latinskt tangentbord.</p>
<p class="p">För att välja en inmatningsmetod, högerklicka på textkomponenten och i menyn <span class="gui">Inmatningsmetod</span> välj inmatningsmetoden du vill använda. Det finns ingen standardinmatningsmetod så läs i dokumentationen för inmatningsmetoder om hur de används.</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="tips.html" title="Tips och tricks">Tips och tricks</a><span class="desc"> — <span class="link"><a href="tips-specialchars.html" title="Mata in speciella tecken">Specialtecken</a></span>, <span class="link"><a href="mouse-middleclick.html" title="Mittenklick">genvägar för mittenklick</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="keyboard-layouts.html" title="Använd alternativa tangentbordslayouter">Använd alternativa tangentbordslayouter</a><span class="desc"> — Lägg till tangentbordslayouter och växla mellan dem.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
