<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ställ in en skrivare</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.04</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="hardware.html" title="Maskinvara och drivrutiner">Hårdvara</a> » <a class="trail" href="printing.html" title="Utskrifter">Utskrifter</a> › <a class="trail" href="printing.html#setup" title="Ställ in en skrivare">Inställningar</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Ställ in en skrivare</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">Du kan ställa in en nätverksansluten eller USB-ansluten skrivare.</p>
<p class="p">För att ställa in en nätverksskrivare:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Skrivaren förutsätts vara ansluten till ditt nätverk. Klicka på ikonen längst till höger i <span class="gui">menylisten</span> och välj <span class="gui">Systeminställningar</span>.</p></li>
<li class="steps"><p class="p">Öppna <span class="gui">Skrivare</span>.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Lägg till</span>.</p></li>
<li class="steps"><p class="p">Om din skrivare finns upptagen i listan över <span class="gui">Enheter</span>, välj den och gå till steg 7.</p></li>
<li class="steps"><p class="p">Du förutsätts veta vilken IP-adress din skrivare har. Välj <span class="gui">Hitta nätverksskrivare</span>, ange IP-adressen i <span class="gui">Host</span>-fältet, och klicka på <span class="gui">Hitta</span>.</p></li>
<li class="steps"><p class="p">Systemet bör nu ha hittat din skrivare. Om inte <span class="gui">Host</span>-fältet visar din IP-adress, ange den igen.</p></li>
<li class="steps"><p class="p">Klicka på <span class="gui">Framåt</span> och vänta medan systemet söker efter drivrutiner.</p></li>
<li class="steps"><p class="p">Välj en drivrutin och installera den.</p></li>
<li class="steps"><p class="p">Du kan anpassa skrivarens namn, beskrivning, och plats om du vill. När du är färdig, klicka på <span class="gui">Verkställ</span>.</p></li>
<li class="steps"><p class="p">Du kan nu skriva ut en testsida eller klicka på <span class="gui">Avbryt</span> för att hoppa över det steget.</p></li>
</ol></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om du har ställt in en nätverksskrivare och den inte vill skriva ut, kontrollera fältet <span class="gui">Enhets-URI</span> i skrivarinställningarna. Det skall visa skrivarens IP-adress. Om inte, korrigera det.</p></div></div></div></div>
<p class="p"> </p>
<p class="p">För att ställa in en USB-ansluten skrivare:</p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">Säkerställ att skrivaren är påslagen.</p></li>
<li class="steps"><p class="p">Anslut skrivaren till ditt system via en lämplig kabel. Det kan förekomma aktivitet på skärmen medan systemet letar efter drivrutiner och du kan bli tillfrågad att autentisera dig för att installera dem.</p></li>
<li class="steps"><p class="p">Ett meddelande kommer visas när systemet har slutfört skrivarinstallationen. Välj <span class="gui">Skriv ut testsida</span> för att skriva ut en testsida, eller <span class="gui">Alternativ</span> för att göra ytterligare ändringar bland skrivarens inställningar.</p></li>
<li class="steps"><p class="p">Du kan dela skrivaren i nätverket, om du vill. Öppna <span class="gui">Skrivare</span>, välj <span class="gui">Server</span> ^ <span class="gui">Inställningar...</span> från menylisten och markera <span class="gui">Publicera utdelade skrivare anslutna till detta system</span>.</p></li>
</ol></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om det finns flera olika drivrutiner tillgängliga för din dator kan du ombes välja en av dem. För att använda den rekommenderade drivrutinen, klicka bara <span class="gui">Framåt</span> på skärmarna för tillverkare och modell.</p></div></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">Om systemet inte kan hitta en drivrutin, försök hitta en på skrivartillverkarens webbplats.</p></div></div></div></div>
<p class="p"> </p>
<p class="p">Efter att du installerat skrivaren, kanske du vill <span class="link"><a href="printing-setup-default-printer.html" title="Ställ in standardskrivaren">ändra din standardskrivare</a></span>.</p>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="printing.html#setup" title="Ställ in en skrivare">Ställ in en skrivare</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
