<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Surfa på nätet</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 17.10</span> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Ubuntu Desktop Guide</a> » <a class="trail" href="getting-started.html" title="Komma igång">Börja med GNOME</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="gs-get-online.html" title="Ansluta till nätet">Föregående</a><a class="nextlinks-next" href="gs-connect-online-accounts.html" title="Ansluta till nätkonton">Nästa</a>
</div>
<div class="hgroup"><h1 class="title"><span class="title">Surfa på nätet</span></h1></div>
<div class="region">
<div class="contents"><div class="steps"><div class="inner"><div class="region"><ol class="steps" start="3">
<li class="steps"><p class="p">Klicka på adressfältet längst upp i webbläsarens fönster och skriv in adressen till den webbplats du vill besöka.</p></li>
<li class="steps">
<p class="p">När en webbplats skrivs in börjar webbläsaren söka efter den bland historik och bokmärken, så du behöver inte komma ihåg den exakta adressen.</p>
<p class="p">Om webbplatsen hittas bland historiken eller bokmärkena kommer en rullgardinslista att visas nedanför adressraden.</p>
</li>
<li class="steps"><p class="p">Från rullgardinslistan kan du snabbt välja en webbplats genom att använda piltangenterna.</p></li>
<li class="steps"><p class="p">Efter att du har valt en webbplats, tryck på <span class="key"><kbd>Retur</kbd></span> för att besöka sidan.</p></li>
</ol></div></div></div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="gs-get-online.html" title="Ansluta till nätet">Föregående</a><a class="nextlinks-next" href="gs-connect-online-accounts.html" title="Ansluta till nätkonton">Nästa</a>
</div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="getting-started.html" title="Komma igång">Börja med GNOME</a><span class="desc"> — Är GNOME nytt för dig? Lär dig hur du använder det.</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-browser.html" title="Webbläsare">Webbläsare</a><span class="desc"> — <span class="link"><a href="net-default-browser.html" title="Ändra vilken webbläsare som öppnar webbplatser som standard">Ändra standardwebbläsare</a></span>, <span class="link"><a href="net-install-flash.html" title="Installera insticksmodulen Flash">installera Flash</a></span>…</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
