<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ljud, video och bilder</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<span style="color: #333">Ubuntu 19.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Ljud, video och bilder</span></h1></div>
<div class="region">
<div class="contents"></div>
<div id="sound" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Grundläggande ljud</span></h2></div>
<div class="region">
<div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="sound-broken.html.sv" title="Ljudproblem"><span class="title">Ljudproblem</span><span class="linkdiv-dash"> — </span><span class="desc">Felsök problem som att inte få ljud eller få dåligt ljudkvalitet.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="sound-usespeakers.html.sv" title="Använd andra högtalar eller hörlurar"><span class="title">Använd andra högtalar eller hörlurar</span><span class="linkdiv-dash"> — </span><span class="desc">Anslut högtalare eller hörlurar och välj en annan standard ljudutmatningsenhet.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="sound-usemic.html.sv" title="Använd en annan mikrofon"><span class="title">Använd en annan mikrofon</span><span class="linkdiv-dash"> — </span><span class="desc">Använd en analog eller USB-mikrofon och välj standardingångsenhet.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="sound-alert.html.sv" title="Välj eller inaktivera larmljudet"><span class="title">Välj eller inaktivera larmljudet</span><span class="linkdiv-dash"> — </span><span class="desc">Välj ett ljud som spelar för meddelanden, ställa in larmljudet eller inaktivera larmljud.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="sound-volume.html.sv" title="Ändra ljudvolymen"><span class="title">Ändra ljudvolymen</span><span class="linkdiv-dash"> — </span><span class="desc">Ställ in ljudvolymen för datorn och kontrollera volymen för varje program.</span></a></div>
</div>
</div></div></div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h3><span class="title">Mer information</span></h3></div>
<div class="region"><ul><li class="links ">
<a href="prefs.html.sv" title="Inställningar för användare och system">Inställningar för användare och system</a><span class="desc"> — <span class="link"><a href="keyboard.html.sv" title="Tangentbord">Tangentbord</a></span>, <span class="link"><a href="mouse.html.sv" title="Mus &amp; styrplatta">mus &amp; styrplatta</a></span>, <span class="link"><a href="prefs-display.html.sv" title="Visning och skärm">visning</a></span>, <span class="link"><a href="prefs-language.html.sv" title="Region &amp; språk">språk</a></span>, <span class="link"><a href="user-accounts.html.sv" title="Användarkonton">användarkonton</a></span>…</span>
</li></ul></div>
</div></div></div>
</div>
</div>
</div></div>
<div id="music" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Musik och bärbara ljudspelare</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="music-cantplay-drm.html.sv" title="Jag kan inte spela låtarna jag köpt från en nätmusikaffär"><span class="title">Jag kan inte spela låtarna jag köpt från en nätmusikaffär</span><span class="linkdiv-dash"> — </span><span class="desc">Stöd för det filformatet kanske inte är installerat eller så kan låtarna vara ”kopieringsskyddade”.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="music-player-ipodtransfer.html.sv" title="Låtar visas inte på min iPod när jag kopierar över dem"><span class="title">Låtar visas inte på min iPod när jag kopierar över dem</span><span class="linkdiv-dash"> — </span><span class="desc">Använd en mediaspelare för att kopiera låtarna och koppla säkert från iPod:en efteråt.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="music-player-newipod.html.sv" title="Min nya iPod fungerar inte"><span class="title">Min nya iPod fungerar inte</span><span class="linkdiv-dash"> — </span><span class="desc">Helt nya iPods måste ställas in via iTunes-programvaran innan du kan använda dem.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="files-autorun.html.sv" title="Öppna program för enheter eller diskar"><span class="title">Öppna program för enheter eller diskar</span><span class="linkdiv-dash"> — </span><span class="desc">Kör automatiskt program för cd och dvd, kameror, musikspelare, och andra enheter och media.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div id="photos" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Foton och digitalkameror</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="hardware-cardreader.html.sv" title="Problem med mediakortsläsare"><span class="title">Problem med mediakortsläsare</span><span class="linkdiv-dash"> — </span><span class="desc">Felsök mediakortsläsare</span></a></div></div>
<div class="links-twocolumn"><div class="linkdiv "><a class="linkdiv" href="files-autorun.html.sv" title="Öppna program för enheter eller diskar"><span class="title">Öppna program för enheter eller diskar</span><span class="linkdiv-dash"> — </span><span class="desc">Kör automatiskt program för cd och dvd, kameror, musikspelare, och andra enheter och media.</span></a></div></div>
</div></div></div></div></div>
</div></div>
<div id="videos" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Videor och videokameror</span></h2></div>
<div class="region"><div class="contents"><div class="links topiclinks"><div class="inner"><div class="region">
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="video-sending.html.sv" title="Andra personer kan inte spela upp videorna jag gjort"><span class="title">Andra personer kan inte spela upp videorna jag gjort</span><span class="linkdiv-dash"> — </span><span class="desc">Kontrollera att de har de korrekta videokodekarna installerade.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="app-cheese.html.sv" title="Skapa roliga bilder och videor med din webbkamera"><span class="title">Skapa roliga bilder och videor med din webbkamera</span><span class="linkdiv-dash"> — </span><span class="desc">Det är lite som ditt privata fotobås.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="video-dvd.html.sv" title="Varför spelas inte dvd-filmer upp?"><span class="title">Varför spelas inte dvd-filmer upp?</span><span class="linkdiv-dash"> — </span><span class="desc">Du kanske inte har rätt kodekar installerade eller så kan dvd:n vara från fel region.</span></a></div>
</div>
<div class="links-twocolumn">
<div class="linkdiv "><a class="linkdiv" href="files-autorun.html.sv" title="Öppna program för enheter eller diskar"><span class="title">Öppna program för enheter eller diskar</span><span class="linkdiv-dash"> — </span><span class="desc">Kör automatiskt program för cd och dvd, kameror, musikspelare, och andra enheter och media.</span></a></div>
<div class="linkdiv "><a class="linkdiv" href="video-dvd-restricted.html.sv" title="Hur aktiverar jag begränsade kodekar för DVD-uppspelning?"><span class="title">Hur aktiverar jag begränsade kodekar för DVD-uppspelning?</span><span class="linkdiv-dash"> — </span><span class="desc">De flesta kommersiella DVD-skivor är krypterade och kommer inte spelas upp utan avkrypteringsprogram.</span></a></div>
</div>
</div></div></div></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="index.html.sv" title="Handbok för Ubuntu-skrivbordet">Handbok för Ubuntu-skrivbordet</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
