<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Varför kopplar mitt trådlösa nätverk ner hela tiden?</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="highlight.pack.js"></script><script>
document.addEventListener('DOMContentLoaded', function() {
  var matches = document.querySelectorAll('code.syntax')
  for (var i = 0; i < matches.length; i++) {
    hljs.highlightBlock(matches[i]);
  }
}, false);</script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><script>
      function englishPageVersion() {

        var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = "index.html.en";
	} else {
		window.location = href.replace(/\.html.*/, ".html.en");
	}
	 return false;
      }

      function browserPreferredLanguage() {
	var href = window.location.href;
	if (href.slice(-1) == "/") {
		window.location = href;
	} else {
		window.location = href.replace(/\.html.*/, ".html");
	}
	return false;
      }
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://canonical.com/partners">Partners</a></li>
<li><a href="https://ubuntu.com/community/support">Support</a></li>
<li><a href="https://ubuntu.com/community">Community</a></li>
<li><a href="https://ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://ubuntu.com/community/contribute">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation">
<div class="trail">
<span style="color: #333">Ubuntu 24.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk</a> » <a class="trail" href="net-problem.html.sv" title="Nätverksproblem">Nätverksproblem</a> » </div>
<div class="trail">
<span style="color: #333">Ubuntu 24.04</span> » <a class="trail" href="index.html.sv" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Hjälp"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="net.html.sv" title="Nätverk, webb &amp; e-post">Nätverk</a> » <a class="trail" href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlösa nätverk</a> » </div>
</div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup pagewide"><h1 class="title"><span class="title">Varför kopplar mitt trådlösa nätverk ner hela tiden?</span></h1></div>
<div class="region">
<div class="contents pagewide"><p class="p">Du kan komma att upptäcka att du har blir frånkopplad från ett trådlöst nätverk även om du ville fortsätta vara ansluten. Din dator kommer normalt att försöka återansluta till nätverket igen så snart detta händer (nätverksikonen i systemraden kommer att visa tre punkter om den försöker återansluta), men det kan vara irriterande, speciellt om du använde internet just då.</p></div>
<section id="signal"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Svag trådlös signal</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">En vanlig orsaka till att man blir frånkopplad från ett trådlöst nätverk är att du har låg signal. Trådlösa nätverk har en begränsad räckvidd, så om du är alltför långt borta från den trådlösa basstationen kanske du inte får tillräckligt stark signal för att upprätthålla en anslutning. Väggar och andra objekt mellan dig och basstationen kan också försvaga signalen.</p>
<p class="p">Nätverksikonen i systemraden visar hur stark din trådlösa signal är. Om signalen ser låg ut, prova att flytta närmare den trådlösa basstationen.</p>
</div></div>
</div></section><section id="network"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Nätverksanslutningen etablerades inte ordentligt</span></h2></div>
<div class="region"><div class="contents pagewide">
<p class="p">Ibland när du ansluter till ett trådlöst nätverk kan det se ut som om du har lyckats ansluta först, men du blir frånkopplad strax efteråt. Detta händer vanligtvis för att din dator bara delvis lyckades ansluta till nätverket — den lyckades etablera en anslutning, men lyckades inte slutföra anslutningen av någon anledning och blev därför frånkopplad.</p>
<p class="p">Ett möjligt skäl till detta är att du skrivit in fel lösenordsfras för det trådlösa nätverket, eller att din dator inte tilläts använda nätverket (till exempel på grund av att nätverket kräver ett användarnamn för att logga in).</p>
</div></div>
</div></section><section id="hardware"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Otillförlitliga trådlös hårdvara/drivrutiner</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">Viss trådlös nätverkshårdvara kan vara lite otillförlitlig. Trådlösa nätverk är komplicerade så trådlösa kort och basstationen stöter ibland på mindre problem och kan tapp anslutningar. Detta är irriterande men händer ganska regelbundet med många enheter. Om du blir frånkopplad från trådlösa nätverk ibland kan detta vara skälet. Om det händer regelbundet bör du överväga att skaffa annan hårdvara.</p></div></div>
</div></section><section id="busy"><div class="inner">
<div class="hgroup pagewide"><h2 class="title"><span class="title">Hektiska trådlösa nätverk</span></h2></div>
<div class="region"><div class="contents pagewide"><p class="p">Trådlösa nätverk på hektiska platser (exempelvis på universitet och caféer) har ofta många datorer som försöker anslut till dem samtidigt. Ibland kan dessa nätverk blir alltför upptagna och kanske inte kan hantera alla de datorer som försöker ansluta, så vissa blir nerkopplade.</p></div></div>
</div></section><section class="links" role="navigation"><div class="inner">
<div class="hgroup pagewide"></div>
<div class="contents pagewide">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul>
<li class="links ">
<a href="net-problem.html.sv" title="Nätverksproblem">Nätverksproblem</a><span class="desc"> — Lös problem med anslutningen till trådlösa och trådbundna nätverk.</span>
</li>
<li class="links ">
<a href="net-wireless.html.sv" title="Trådlösa nätverk">Trådlösa nätverk</a><span class="desc"> — Anslut till trådlösa nätverk, inklusive dolda nätverk och nätverk består av en surfzon från en telefon.</span>
</li>
</ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="net-wireless-connect.html.sv" title="Anslut till ett trådlöst nätverk">Anslut till ett trådlöst nätverk</a><span class="desc"> — Nå internet — trådlöst.</span>
</li></ul></div>
</div></div>
</div>
</div></section>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer">
<p style="padding-bottom: 0.4em">You can choose the <b>displayed language</b> by adding a language suffix to the web address so it ends with e.g. <tt>.html.en</tt> or <tt>.html.de</tt>.<br>
          If the web address has no language suffix, the preferred language specified in your web browser's settings is used. For your convenience:<br>

          [ <a title="English page version" href="#" onClick="englishPageVersion();">Change to English Language</a> | 
          <a title="Language selected by browser" href="#" onClick="browserPreferredLanguage()">Change to Browser's Preferred Language</a> ]</p>
<p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p>
</div>
</div>
</body>
</html>
