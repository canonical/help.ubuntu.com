<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Skriv speciella tecken</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="tips.html" title="Tips och tricks">Tips och tricks</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">Skriv speciella tecken</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">You can enter and view thousands of characters from most of the 
  world's writing systems, even those not found on your keyboard. This 
  page lists some different ways you can enter special characters.</p>
<div role="navigation" class="links sectionlinks"><div class="inner">
<div class="title title-links"><h2><span class="title">Methods to enter characters</span></h2></div>
<div class="region"><ul>
<li class="links "><a href="tips-specialchars.html#charmap" title="Character map">Character map</a></li>
<li class="links "><a href="tips-specialchars.html#ctrlshiftu" title="Code points">Code points</a></li>
<li class="links "><a href="tips-specialchars.html#sources" title="Input sources">Input sources</a></li>
</ul></div>
</div></div>
</div>
<div id="charmap" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Character map</span></h2></div>
<div class="region"><div class="contents">
<p class="p">GNOME comes with a character map application that allows you to 
    browse all the characters in Unicode. Use the character map to find 
    the character you want, and then copy and paste it to wherever you 
    need it.</p>
<p class="p">You can find <span class="app">Character Map</span> in the <span class="gui">Dash</span>.
    For more information on the character map, see the
    <span class="link"><a href="https://help.gnome.org/users/gucharmap/stable/" title="https://help.gnome.org/users/gucharmap/stable/">Character Map Manual</a></span>.</p>
</div></div>
</div></div>
<div id="ctrlshiftu" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Code points</span></h2></div>
<div class="region"><div class="contents">
<p class="p">You can enter any Unicode character using only your keyboard with 
    the numeric code point of the character. Every character is identified 
    by a four-character code point. To find the code point for a 
    character, find the character in the character map application and 
    look in the status bar or the <span class="gui">Character Details</span> tab. The 
    code point is the four characters after <span class="gui">U+</span>.</p>
<p class="p">To enter a character by its code point, hold down <span class="key"><kbd>Ctrl</kbd></span> 
    and <span class="key"><kbd>Shift</kbd></span>, type <span class="key"><kbd>u</kbd></span> followed by the four-character 
    code point, then release <span class="key"><kbd>Ctrl</kbd></span> and <span class="key"><kbd>Shift</kbd></span>. If you 
    often use characters that you can't easily access with other methods, 
    you might find it useful to memorize the code point for those 
    characters so you can enter them quickly.</p>
</div></div>
</div></div>
<div id="sources" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Input sources</span></h2></div>
<div class="region"><div class="contents"><p class="p">You can make your keyboard behave like the keyboard for another 
    language, regardless of the letters printed on the keys. You can even 
    switch between different input sources using an icon in the menu 
    bar. To learn how, see <span class="link"><a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">Använd alternativa inmatningskällor</a></span>.</p></div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents">
<div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="tips.html" title="Tips och tricks">Tips och tricks</a><span class="desc"> — <span class="link"><a href="tips-specialchars.html" title="Skriv speciella tecken">Speciella tecken</a></span>, <span class="link"><a href="mouse-middleclick.html" title="Mittenklick">mittenklick</a></span>…</span>
</li></ul></div>
</div></div>
<div class="links seealsolinks"><div class="inner">
<div class="title"><h2><span class="title">Se även</span></h2></div>
<div class="region"><ul><li class="links ">
<a href="keyboard-layouts.html" title="Använd alternativa inmatningskällor">Använd alternativa inmatningskällor</a><span class="desc"> — Lägg till indatakällor och växla mellan dem.</span>
</li></ul></div>
</div></div>
</div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
