<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Manager</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="https://partners.ubuntu.com">Partners</a></li>
<li><a href="https://www.ubuntu.com/support/community-support">Support</a></li>
<li><a href="https://community.ubuntu.com">Community</a></li>
<li><a href="https://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="https://community.ubuntu.com/t/contribute/26">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../16.04" class="trail">Ubuntu 16.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="cgroups.html" title="Control Groups">Control Groups</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups-delegation.html" title="Delegation">Föregående</a><a class="nextlinks-next" href="cgroups-resources.html" title="Resurser">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Manager</h1></div>
<div class="region"><div class="contents">
<p class="para">
The cgroup manager (cgmanager) provides a D-Bus service allowing
programs and users to administer cgroups without needing direct
knowledge of or access to the cgroup filesystem.  For requests
from tasks in the same namespaces as the manager, the manager can
directly perform the needed security checks to ensure that requests
are legitimate.  For other requests - such as those from a task in
a container - enhanced D-Bus requests must be made, where process-,
user- and group-ids are passed as SCM_CREDENTIALS, so that the kernel
maps the identifiers to their global host values.
  </p>
<p class="para">
To fascilitate the use of simple D-Bus calls from all users, a
'cgroup manager proxy' (cgproxy) is automatically started when in
a container.  The proxy accepts standard D-Bus requests from tasks
in the same namespaces as itself, and converts them to 
SCM-enhanced D-Bus requests which it passes on to the cgmanager.
  </p>
<p class="para">
A simple example of creating a new cgroup in which to run a
cpu-intensive compile would look like:
  </p>
<div class="screen"><pre class="contents "><span class="cmd command">
cgm create cpuset build1
cgm movepid cpuset build1 $$
cgm setvalue cpuset build1 cpuset.cpus 1
make
</span></pre></div>
</div></div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="cgroups-delegation.html" title="Delegation">Föregående</a><a class="nextlinks-next" href="cgroups-resources.html" title="Resurser">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
