<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>Ubuntu Cloud</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Ubuntu serverguide">Ubuntu serverguide</a> » <a class="trail" href="virtualization.html" title="Virtualisering">Virtualisering</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="links nextlinks">
<a class="nextlinks-prev" href="cloud-images-and-uvtool.html" title="Cloud images and uvtool">Föregående</a><a class="nextlinks-next" href="lxc.html" title="LXC">Nästa</a>
</div>
<div class="hgroup"><h1 class="title">Ubuntu Cloud</h1></div>
<div class="region">
<div class="contents"><p class="para"><span class="app application">Cloud computing</span> is a computing model that
    allows vast pools of resources to be allocated on-demand. These resources
    such as storage, computing power, network and software are abstracted and
    delivered as a service over the Internet anywhere, anytime. These services
    are billed per time consumed similar to the ones used by public services
    such as electricity, water and telephony. <span class="app application">Ubuntu Cloud
    Infrastructure</span> uses OpenStack open source software to help
    build highly scalable, cloud computing for both public and private
    clouds.</p></div>
<div class="links sectionlinks" role="navigation"><ul>
<li class="links"><a class="xref" href="ubuntucloud.html#ubuntu-cloud-installation" title="Installation and Configuration">Installation and Configuration</a></li>
<li class="links"><a class="xref" href="ubuntucloud.html#ubuntu-cloud-troubleshooting" title="Support and Troubleshooting">Support and Troubleshooting</a></li>
<li class="links"><a class="xref" href="ubuntucloud.html#ubuntu-cloud-resources" title="Resurser">Resurser</a></li>
</ul></div>
<div class="sect2 sect" id="ubuntu-cloud-installation"><div class="inner">
<div class="hgroup"><h2 class="title">Installation and Configuration</h2></div>
<div class="region"><div class="contents"><p class="para">
	    Due to the current high rate of development of this complex technology
	    we refer the reader to <a href="http://docs.openstack.org/havana/install-guide/install/apt/content/" class="ulink" title="http://docs.openstack.org/havana/install-guide/install/apt/content/">
	    upstream documentation</a> for all matters concerning installation and configuration.
    </p></div></div>
</div></div>
<div class="sect2 sect" id="ubuntu-cloud-troubleshooting"><div class="inner">
<div class="hgroup"><h2 class="title">Support and Troubleshooting</h2></div>
<div class="region"><div class="contents">
<p class="para">Community Support</p>
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
          <p class="para"><a href="https://launchpad.net/~openstack" class="ulink" title="https://launchpad.net/~openstack">OpenStack
          Mailing list</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para"><a href="http://wiki.openstack.org" class="ulink" title="http://wiki.openstack.org">The OpenStack Wiki
          search</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para"><a href="https://bugs.launchpad.net/nova" class="ulink" title="https://bugs.launchpad.net/nova">Launchpad bugs
          area</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para">Join the IRC channel #openstack on freenode.</p>
        </li>
</ul></div>
</div></div>
</div></div>
<div class="sect2 sect" id="ubuntu-cloud-resources"><div class="inner">
<div class="hgroup"><h2 class="title">Resurser</h2></div>
<div class="region"><div class="contents">
<div class="list itemizedlist"><ul class="list itemizedlist">
<li class="list itemizedlist">
          <p class="para"><a href="http://en.wikipedia.org/wiki/Cloud_computing#Service_Models" class="ulink" title="http://en.wikipedia.org/wiki/Cloud_computing#Service_Models">Cloud
          Computing - Service models</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para"><a href="http://www.openstack.org/software/openstack-compute/" class="ulink" title="http://www.openstack.org/software/openstack-compute/">OpenStack
          Compute</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para"><a href="http://docs.openstack.org/diablo/openstack-compute/starter/content/GlanceMS-d2s21.html" class="ulink" title="http://docs.openstack.org/diablo/openstack-compute/starter/content/GlanceMS-d2s21.html">OpenStack
          Image Service</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para"><a href="http://docs.openstack.org/trunk/openstack-object-storage/admin/content/index.html" class="ulink" title="http://docs.openstack.org/trunk/openstack-object-storage/admin/content/index.html">OpenStack Object
          Storage Administration Guide</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para"><a href="http://docs.openstack.org/trunk/openstack-object-storage/admin/content/installing-openstack-object-storage-on-ubuntu.html" class="ulink" title="http://docs.openstack.org/trunk/openstack-object-storage/admin/content/installing-openstack-object-storage-on-ubuntu.html">Installing
          OpenStack Object Storage on Ubuntu</a></p>
        </li>
<li class="list itemizedlist">
          <p class="para"><a href="http://cloudglossary.com/" class="ulink" title="http://cloudglossary.com/">http://cloudglossary.com/</a></p>
        </li>
</ul></div>
<p class="para"></p>
</div></div>
</div></div>
</div>
<div class="links nextlinks">
<a class="nextlinks-prev" href="cloud-images-and-uvtool.html" title="Cloud images and uvtool">Föregående</a><a class="nextlinks-next" href="lxc.html" title="LXC">Nästa</a>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this serverguide documentation, <a href="https://bugs.launchpad.net/serverguide">file a bug report</a>.</p></div>
</div>
</body>
</html>
