<!DOCTYPE html>
<html lang=sv>
<head>
<meta http-equiv="Content-Type" content="text/html; charset=UTF-8">
<title>I forgot my password!</title>
<link rel="stylesheet" type="text/css" href="sv.css">
<script type="text/javascript" src="jquery.js"></script><script type="text/javascript" src="jquery.syntax.js"></script><script type="text/javascript" src="yelp.js"></script>
</head>
<body id="home">
<script src="https://ssl.google-analytics.com/urchin.js" type="text/javascript"></script><script type="text/javascript">
        _uacct = "UA-1018242-8";
        urchinTracker();
      </script><div id="container">
<div id="container-inner">
<div id="mothership"><ul>
<li><a href="http://www.ubuntu.com/partners">Partners</a></li>
<li><a href="http://www.ubuntu.com/support">Support</a></li>
<li><a href="http://www.ubuntu.com/community">Community</a></li>
<li><a href="http://www.ubuntu.com">Ubuntu.com</a></li>
</ul></div>
<div id="header">
<h1 id="ubuntu-header"><a href="https://help.ubuntu.com/">Ubuntu Documentation</a></h1>
<ul id="main-menu">
<li><a class="main-menu-item current" href="../../">Official Documentation</a></li>
<li><a href="https://help.ubuntu.com/community/CommunityHelpWiki">Community Help Wiki</a></li>
<li><a href="http://community.ubuntu.com/contribute/documentation/">Contribute</a></li>
</ul>
</div>
<div id="menu-search"><div id="search-box">
<noscript><form action="https://www.google.com/cse" id="cse-search-box"><div>
<input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq"><input type="hidden" name="ie" value="UTF-8"><input type="text" name="q" size="21"><input type="submit" name="sa" value="Search">
</div></form></noscript>
<script>
                document.write('<form action="../../search.html" id="cse-search-box">');
                document.write('  <div>');
                document.write('    <input type="hidden" name="cof" value="FORID:9">');
                document.write('    <input type="hidden" name="cx" value="003883529982892832976:e2vwumte3fq">');
                document.write('    <input type="hidden" name="ie" value="UTF-8">');
                document.write('    <input type="text" name="q" size="21">');
                document.write('    <input type="submit" name="sa" value="Search">');
                document.write('  </div>');
                document.write('</form>');
              </script>
</div></div>
<div class="trails" role="navigation"><div class="trail">
<a href="../../14.04" class="trail">Ubuntu 14.04</a> » <a class="trail" href="index.html" title="Handbok för Ubuntu-skrivbordet"><span class="media"><span class="media media-image"><img src="figures/ubuntu-logo.png" height="16" width="16" class="media media-inline" alt="Help"></span></span> Handbok för Ubuntu-skrivbordet</a> » <a class="trail" href="prefs.html" title="Inställningar för användare och system">Settings</a> » <a class="trail" href="user-accounts.html" title="Användarkonton">Users</a> › <a class="trail" href="user-accounts.html#passwords" title="Lösenord">Lösenord</a> » </div></div>
<div id="cwt-content" class="clearfix content-area"><div id="page">
<div id="content">
<div class="hgroup"><h1 class="title"><span class="title">I forgot my password!</span></h1></div>
<div class="region">
<div class="contents">
<p class="p">
     It is important to choose not only <span class="link"><a href="user-goodpassword.html" title="Välj ett säkert lösenord">a good
 and secure password</a></span>, but also one that you can remember. If you have
 forgotten the password to log in to your computer account, you can follow the
 following steps to reset it.
  </p>
<div class="note note-important" title="Viktigt"><div class="inner"><div class="region"><div class="contents"><p class="p">
     If you have an encrypted home directory, you will not be able to reset a
 forgotten password.
  </p></div></div></div></div>
<p class="p">
  If you simply want to change your password, see <span class="link"><a href="user-changepassword.html" title="Välj ditt lösenord">Välj ditt lösenord</a></span>.
  </p>
<div role="navigation" class="links sectionlinks"><div class="inner"><div class="region"><ul>
<li class="links "><a href="user-forgottenpassword.html#reset-password-grub2" title="Reset password using Grub">Reset password using Grub</a></li>
<li class="links "><a href="user-forgottenpassword.html#live-cd" title="Reset password using a Live CD or USB">Reset password using a Live CD or USB</a></li>
<li class="links "><a href="user-forgottenpassword.html#delete-keyring" title="Get rid of the keyring">Get rid of the keyring</a></li>
</ul></div></div></div>
</div>
<div id="reset-password-grub2" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Reset password using Grub</span></h2></div>
<div class="region"><div class="contents">
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps">
<p class="p">
           Restart your computer, and hold down <span class="key"><kbd>Shift</kbd></span> during bootup
 to get into the Grub menu.
           </p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">
           If you have a dual-boot machine and you choose at boot time which
 operating system to boot into, the Grub menu should appear without the need to
 hold down <span class="key"><kbd>Shift</kbd></span>.
           </p></div></div></div></div>
<div class="note" title="Anteckning"><div class="inner"><div class="region"><div class="contents"><p class="p">If you are unable to get into the Grub boot menu, and therefore cannot choose to boot into recovery mode, you can <span class="link"><a href="user-forgottenpassword.html#live-cd" title="Reset password using a Live CD or USB">use a live CD to reset your user password</a></span>.
           </p></div></div></div></div>
</li>
<li class="steps"><p class="p">
           Press the down arrow on your keyboard to highlight the line that ends with the words 'recovery mode',
then press <span class="key"><kbd>Enter</kbd></span>.
           </p></li>
<li class="steps"><p class="p">
           Your computer will now begin the boot process. After a few moments, a <span class="gui">Recovery Menu</span> will appear.
           Use your down arrow key to highlight <span class="gui">root</span> and press <span class="key"><kbd>Enter</kbd></span>.
           </p></li>
<li class="steps">
<p class="p">
           At the <span class="cmd">#</span> symbol, type:
           </p>
<p class="p">
           <span class="cmd">passwd <span class="var">username</span></span>, where <span class="var">username</span> is the username of the account you're changing the password for.
           </p>
</li>
<li class="steps"><p class="p">
           You will be prompted to enter a new UNIX password, and to confirm the new password.
           </p></li>
<li class="steps">
<p class="p">
           Then type:
           </p>
<p class="p">
           # <span class="cmd">reboot</span>
           </p>
</li>
</ol></div></div></div>
<p class="p">
       After you successfully log in, you will not be able to access your keyring
 (since you don't remember the old password).  This means that all your saved
 passwords for wireless networks, jabber accounts, etc. will no longer be
 accessible.  You will need to <span class="link"><a href="#delete-keyring" title="Get rid of the keyring">delete the old
 keyring</a></span> and start a new one.
     </p>
</div></div>
</div></div>
<div id="live-cd" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Reset password using a Live CD or USB</span></h2></div>
<div class="region"><div class="contents">
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">
           Boot the Live CD or USB.
           </p></li>
<li class="steps"><p class="p">Montera din enhet.</p></li>
<li class="steps"><p class="p">
           Press <span class="keyseq"><span class="key"><kbd>Alt</kbd></span>+<span class="key"><kbd>F2</kbd></span></span> to get the <span class="gui">Run
           Application</span> window.
           </p></li>
<li class="steps">
<p class="p">
           Type <span class="cmd">gksu nautilus</span> to launch the file manager with system-wide privileges.
           </p>
<div class="note note-tip" title="Tips"><div class="inner"><div class="region"><div class="contents"><p class="p">
             Within the drive you just mounted, you can check that it is the right
             drive by clicking <span class="gui"> home </span> and then your username.
           </p></div></div></div></div>
</li>
<li class="steps">
<p class="p">
           Go to the top-level directory of the mounted drive.  Then go into the <span class="gui">etc</span> directory.
           </p>
<p class="p">
           Locate the 'shadow' file and make a backup copy:
           </p>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">
           Right-click on the shadow file and select <span class="gui">copy</span>.
           </p></li>
<li class="steps"><p class="p">
            Then right-click in the empty space and select <span class="gui">paste</span>.
           </p></li>
<li class="steps"><p class="p">
                      <span class="link"><a href="files-rename.html" title="Byt namn på en fil eller mapp">Rename</a></span> the backup "shadow.bak".
           </p></li>
</ol></div></div></div>
</li>
<li class="steps"><p class="p">
           Edit the original "shadow" file with a text editor.
           </p></li>
<li class="steps">
<p class="p">
           Find your username for which you have forgotten the password.  It
 should look something like this (the characters after the colon will be different):
           </p>
<p class="p">
           username:$1$2abCd0E or
           </p>
<p class="p">
           username:$1$2abCd0E:13721a:0:99999:7:::
           </p>
</li>
<li class="steps">
<p class="p">
         Delete the characters after the first colon and before the second
 colon. This will remove the password for the account.
           </p>
<p class="p">
           Save the file, exit out of everything and reboot your computer without
 the live CD or USB.
           </p>
</li>
<li class="steps"><p class="p">
           When you boot back into your installation, click your name in the menu bar. Open <span class="gui">My Account</span> and reset your password.
           </p></li>
<li class="steps"><p class="p">
            For <span class="gui">Current password</span> do not enter anything, as your
 current password is blank.  Just click <span class="gui">Authenticate</span> and enter a new
 password.
          </p></li>
</ol></div></div></div>
<p class="p">
       After you successfully log in, you will not be able to access your keyring
 (since you don't remember the old password).  This means that all your saved
 passwords for wireless networks, jabber accounts, etc. will no longer be
 accessible.  You will need to <span class="link"><a href="#delete-keyring" title="Get rid of the keyring">delete the old
 keyring</a></span> and start a new one.
     </p>
</div></div>
</div></div>
<div id="delete-keyring" class="sect"><div class="inner">
<div class="hgroup"><h2 class="title"><span class="title">Get rid of the keyring</span></h2></div>
<div class="region"><div class="contents">
<div class="note note-warning" title="Varning"><div class="inner"><div class="region"><div class="contents"><p class="p">This will delete all your saved passwords for wireless
    networks, instant messaging accounts, etc. Only do this if you can't remember
    the password you used for your keyring.</p></div></div></div></div>
<div class="steps"><div class="inner"><div class="region"><ol class="steps">
<li class="steps"><p class="p">
    Go to your Home folder by typing 'home' in the <span class="gui">Dash</span>.
   </p></li>
<li class="steps"><p class="p">
    Press <span class="keyseq"><span class="key"><kbd>Ctrl</kbd></span>+<span class="key"><kbd>h</kbd></span></span> (or click
 <span class="guiseq"><span class="gui">View</span> ▸ <span class="gui">Show Hidden Files</span></span>.)
   </p></li>
<li class="steps"><p class="p">
    Double click on the folder <span class="file">~/.local/share</span>.
   </p></li>
<li class="steps"><p class="p">
   Double click on the folder called keyrings.
   </p></li>
<li class="steps"><p class="p">
   Delete any files you find in the keyrings folder.
   </p></li>
<li class="steps"><p class="p">Starta om datorn.</p></li>
</ol></div></div></div>
<p class="p">
 After you restart and log in you will be asked to enter your wireless networks
 password.
</p>
</div></div>
</div></div>
<div class="sect sect-links" role="navigation">
<div class="hgroup"></div>
<div class="contents"><div class="links guidelinks"><div class="inner">
<div class="title"><h2><span class="title">Mer information</span></h2></div>
<div class="region"><ul><li class="links "><a href="user-accounts.html#passwords" title="Lösenord">Lösenord</a></li></ul></div>
</div></div></div>
</div>
</div>
<div class="clear"></div>
</div>
<div id="pagebottom"></div>
</div></div>
</div>
<div id="footer"><p>The material in this document is available under a free license, see <a href="../../legal.html">Legal</a> for details.<br>
          For information on contributing see the <a href="https://wiki.ubuntu.com/DocumentationTeam">Ubuntu Documentation Team wiki page</a>.
          To report errors in this documentation, <a href="https://bugs.launchpad.net/ubuntu/+source/ubuntu-docs">file a bug</a>.</p></div>
</div>
</body>
</html>
